magic
tech scmos
timestamp 1497186066
<< nwell >>
rect 0 36 99 75
<< pwell >>
rect 0 -3 99 36
<< ntransistor >>
rect 20 21 22 29
rect 36 21 38 25
rect 44 21 46 25
rect 52 21 54 25
rect 62 21 64 25
rect 78 21 80 29
<< ptransistor >>
rect 20 43 22 59
rect 36 55 38 59
rect 44 55 46 59
rect 52 55 54 59
rect 62 55 64 59
rect 78 43 80 59
<< ndiffusion >>
rect 15 27 20 29
rect 19 23 20 27
rect 15 21 20 23
rect 22 25 27 29
rect 73 25 78 29
rect 22 21 23 25
rect 35 21 36 25
rect 38 21 39 25
rect 43 21 44 25
rect 46 21 47 25
rect 51 21 52 25
rect 54 21 57 25
rect 61 21 62 25
rect 64 21 65 25
rect 77 21 78 25
rect 80 27 85 29
rect 80 23 81 27
rect 80 21 85 23
<< pdiffusion >>
rect 15 58 20 59
rect 19 44 20 58
rect 15 43 20 44
rect 22 55 23 59
rect 35 55 36 59
rect 38 55 39 59
rect 43 55 44 59
rect 46 55 47 59
rect 51 55 52 59
rect 54 55 57 59
rect 61 55 62 59
rect 64 55 65 59
rect 77 55 78 59
rect 22 43 27 55
rect 73 43 78 55
rect 80 58 85 59
rect 80 44 81 58
rect 80 43 85 44
<< ndcontact >>
rect 15 23 19 27
rect 23 21 27 25
rect 31 21 35 25
rect 39 21 43 25
rect 47 21 51 25
rect 57 21 61 25
rect 65 21 69 25
rect 73 21 77 25
rect 81 23 85 27
<< pdcontact >>
rect 15 44 19 58
rect 23 55 27 59
rect 31 55 35 59
rect 39 55 43 59
rect 47 55 51 59
rect 57 55 61 59
rect 65 55 69 59
rect 73 55 77 59
rect 81 44 85 58
<< psubstratepcontact >>
rect 23 13 27 17
rect 31 13 35 17
rect 65 13 69 17
rect 73 13 77 17
rect 23 5 27 9
rect 31 5 35 9
rect 65 5 69 9
rect 73 5 77 9
<< nsubstratencontact >>
rect 23 63 27 67
rect 39 63 43 67
rect 47 63 51 67
rect 57 63 61 67
rect 73 63 77 67
<< polysilicon >>
rect 20 59 22 61
rect 36 59 38 61
rect 44 59 46 61
rect 52 59 54 61
rect 62 59 64 61
rect 78 59 80 61
rect 20 39 22 43
rect 36 39 38 55
rect 44 52 46 55
rect 20 29 22 35
rect 36 25 38 35
rect 44 25 46 48
rect 52 39 54 55
rect 52 25 54 35
rect 62 25 64 55
rect 78 29 80 43
rect 20 19 22 21
rect 36 19 38 21
rect 44 19 46 21
rect 52 19 54 21
rect 62 19 64 21
rect 78 19 80 21
<< polycontact >>
rect 42 48 46 52
rect 18 35 22 39
rect 34 35 38 39
rect 52 35 56 39
rect 64 48 68 52
rect 80 35 84 39
<< metal1 >>
rect 1 69 99 75
rect 15 58 19 69
rect 23 67 27 69
rect 39 67 43 69
rect 31 59 35 62
rect 8 39 12 49
rect 15 43 19 44
rect 47 67 51 69
rect 57 67 61 69
rect 73 67 77 69
rect 39 59 43 63
rect 65 59 69 62
rect 23 52 27 55
rect 57 52 61 55
rect 73 52 77 55
rect 23 49 42 52
rect 23 47 27 49
rect 68 48 77 52
rect 73 47 77 48
rect 35 42 65 45
rect 81 58 85 69
rect 81 43 85 44
rect 8 35 18 39
rect 22 35 34 39
rect 56 35 80 38
rect 84 35 89 39
rect 15 27 19 29
rect 15 3 19 23
rect 23 25 27 28
rect 51 28 57 32
rect 47 25 51 28
rect 73 25 77 28
rect 31 17 35 21
rect 23 9 27 13
rect 23 3 27 5
rect 39 18 43 21
rect 57 18 61 21
rect 39 14 61 18
rect 81 27 85 29
rect 65 17 69 21
rect 31 9 35 13
rect 31 3 35 5
rect 65 9 69 13
rect 65 3 69 5
rect 73 9 77 13
rect 73 3 77 5
rect 81 3 85 23
rect 1 -3 99 3
<< m2contact >>
rect 31 62 35 66
rect 8 49 12 53
rect 65 62 69 66
rect 57 48 61 52
rect 23 43 27 47
rect 31 42 35 46
rect 65 41 69 45
rect 73 43 77 47
rect 89 35 93 39
rect 23 28 27 32
rect 47 28 51 32
rect 57 28 61 32
rect 73 28 77 32
<< metal2 >>
rect 7 53 13 54
rect 7 49 8 53
rect 12 49 13 53
rect 7 48 13 49
rect 23 32 27 43
rect 31 46 35 62
rect 46 32 52 33
rect 46 28 47 32
rect 51 28 52 32
rect 57 32 61 48
rect 65 45 69 62
rect 73 32 77 43
rect 88 39 94 40
rect 88 35 89 39
rect 93 35 94 39
rect 88 34 94 35
rect 46 27 52 28
<< m3p >>
rect 2 0 98 72
<< labels >>
rlabel metal1 7 3 7 3 4 gnd
rlabel metal1 7 75 7 75 4 vdd
rlabel metal2 7 48 7 48 1 a
rlabel metal2 88 34 88 34 1 b
rlabel metal2 46 27 46 27 1 out
<< end >>
