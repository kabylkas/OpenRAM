MACRO ecc
    CLASS RING ;
    ORIGIN 66.9 0.0 ;
    FOREIGN  sram 0.0 0.0 ;
    SIZE 232.5 BY 459.3 ;
    SYMMETRY X Y R90 ;
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        SHAPE ABUTMENT ; 
        PORT             
        Layer metal1 ; 
        RECT  0.0 0.0 9.0 459.3 ;
        RECT  157.2 0.0 166.2 459.3 ;
        END             
    END vdd 
    PIN gnd 
        DIRECTION INOUT ; 
        USE GROUND ; 
        SHAPE ABUTMENT ; 
        PORT             
        Layer metal2 ; 
        RECT  95.1 0.0 104.1 459.3 ;
        END             
    END gnd 
    PIN DATA[0] 
        DIRECTION INOUT ; 
        PORT             
        Layer metal3 ; 
        RECT  128.25 0.0 129.75 30.15 ;
        RECT  128.25 0.0 130.05 1.8 ;
        END             
    END DATA[0] 
    PIN DATA[1] 
        DIRECTION INOUT ; 
        PORT             
        Layer metal3 ; 
        RECT  138.45 0.0 139.95 30.15 ;
        RECT  138.45 0.0 140.25 1.8 ;
        END             
    END DATA[1] 
    PIN DATA[2] 
        DIRECTION INOUT ; 
        PORT             
        Layer metal3 ; 
        RECT  148.65 0.0 150.15 30.15 ;
        RECT  148.65 0.0 150.45 1.8 ;
        END             
    END DATA[2] 
    PIN ADDR[0] 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  0.0 73.95 17.1 75.45 ;
        END             
    END ADDR[0] 
    PIN ADDR[1] 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  0.0 63.75 17.1 65.25 ;
        END             
    END ADDR[1] 
    PIN ADDR[2] 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  0.0 53.55 17.1 55.05 ;
        END             
    END ADDR[2] 
    PIN ADDR[3] 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  0.0 43.35 17.1 44.85 ;
        END             
    END ADDR[3] 
    PIN CSb 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  -62.1 86.4 -60.3 88.2 ;
        END             
    END CSb 
    PIN OEb 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  -41.7 86.4 -39.9 88.2 ;
        END             
    END OEb 
    PIN WEb 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  -51.9 86.4 -50.1 88.2 ;
        END             
    END WEb 
    PIN clk 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  -27.15 85.5 105.9 87.0 ;
        RECT  -27.6 85.5 -25.8 87.3 ;
        END             
    END clk 
    OBS 
        Layer  metal1 ; 
        RECT  -10.2 292.65 0.0 293.55 ;
        RECT  157.2 0.0 166.2 459.3 ;
        RECT  0.0 0.0 9.0 459.3 ;
        RECT  51.0 206.4 51.9 209.7 ;
        RECT  51.0 219.9 51.9 223.2 ;
        RECT  51.0 235.8 51.9 239.1 ;
        RECT  51.0 249.3 51.9 252.6 ;
        RECT  51.0 265.2 51.9 268.5 ;
        RECT  51.0 278.7 51.9 282.0 ;
        RECT  51.0 294.6 51.9 297.9 ;
        RECT  51.0 308.1 51.9 311.4 ;
        RECT  51.0 324.0 51.9 327.3 ;
        RECT  51.0 337.5 51.9 340.8 ;
        RECT  51.0 353.4 51.9 356.7 ;
        RECT  51.0 366.9 51.9 370.2 ;
        RECT  51.0 382.8 51.9 386.1 ;
        RECT  51.0 396.3 51.9 399.6 ;
        RECT  51.0 412.2 51.9 415.5 ;
        RECT  51.0 425.7 51.9 429.0 ;
        RECT  88.5 214.35 123.9 215.25 ;
        RECT  88.5 243.75 123.9 244.65 ;
        RECT  88.5 273.15 123.9 274.05 ;
        RECT  88.5 302.55 123.9 303.45 ;
        RECT  88.5 331.95 123.9 332.85 ;
        RECT  88.5 361.35 123.9 362.25 ;
        RECT  88.5 390.75 123.9 391.65 ;
        RECT  88.5 420.15 123.9 421.05 ;
        RECT  74.4 88.8 91.5 89.7 ;
        RECT  74.4 104.7 88.8 105.6 ;
        RECT  74.4 147.6 86.1 148.5 ;
        RECT  74.4 163.5 83.4 164.4 ;
        RECT  114.0 33.3 129.0 34.2 ;
        RECT  108.6 28.65 129.3 29.55 ;
        RECT  111.3 26.25 129.3 27.15 ;
        RECT  114.0 446.4 123.9 447.3 ;
        RECT  116.7 97.95 123.9 98.85 ;
        RECT  119.4 196.05 123.9 196.95 ;
        RECT  123.9 213.75 157.2 214.65 ;
        RECT  123.9 243.15 157.2 244.05 ;
        RECT  123.9 272.55 157.2 273.45 ;
        RECT  123.9 301.95 157.2 302.85 ;
        RECT  123.9 331.35 157.2 332.25 ;
        RECT  123.9 360.75 157.2 361.65 ;
        RECT  123.9 390.15 157.2 391.05 ;
        RECT  123.9 419.55 157.2 420.45 ;
        RECT  123.9 458.4 157.2 459.3 ;
        RECT  123.9 168.75 157.2 169.65 ;
        RECT  123.9 100.05 157.2 100.95 ;
        RECT  123.9 87.3 157.2 88.2 ;
        RECT  129.3 10.35 157.2 11.25 ;
        RECT  138.9 10.35 157.2 11.25 ;
        RECT  149.7 10.35 157.2 11.25 ;
        RECT  0.0 214.35 29.4 215.25 ;
        RECT  0.0 243.75 29.4 244.65 ;
        RECT  0.0 273.15 29.4 274.05 ;
        RECT  0.0 302.55 29.4 303.45 ;
        RECT  0.0 331.95 29.4 332.85 ;
        RECT  0.0 361.35 29.4 362.25 ;
        RECT  0.0 390.75 29.4 391.65 ;
        RECT  0.0 420.15 29.4 421.05 ;
        RECT  0.0 126.15 29.4 127.05 ;
        RECT  0.0 184.95 29.4 185.85 ;
        RECT  95.1 437.1 154.5 438.0 ;
        RECT  101.7 8.1 154.5 9.0 ;
        RECT  29.4 140.85 95.1 141.75 ;
        RECT  29.4 199.65 95.1 200.55 ;
        RECT  75.3 69.15 95.1 70.05 ;
        RECT  75.3 69.15 95.1 70.05 ;
        RECT  75.3 48.75 95.1 49.65 ;
        RECT  75.3 48.75 95.1 49.65 ;
        RECT  123.3 213.6 134.7 214.8 ;
        RECT  124.5 211.5 125.7 213.6 ;
        RECT  127.5 211.5 128.7 212.7 ;
        RECT  130.5 211.5 131.7 212.7 ;
        RECT  133.5 211.5 134.7 213.6 ;
        RECT  127.2 210.6 128.4 211.5 ;
        RECT  124.5 204.9 125.7 210.6 ;
        RECT  127.2 209.4 129.6 210.6 ;
        RECT  127.2 206.1 128.4 209.4 ;
        RECT  130.8 207.9 132.0 211.5 ;
        RECT  130.2 206.7 132.0 207.9 ;
        RECT  130.8 206.1 132.0 206.7 ;
        RECT  126.9 204.9 128.1 206.1 ;
        RECT  131.1 204.9 132.3 206.1 ;
        RECT  133.5 204.9 134.7 210.6 ;
        RECT  129.0 203.4 130.2 203.7 ;
        RECT  123.3 202.2 134.7 203.4 ;
        RECT  125.4 200.1 128.1 201.3 ;
        RECT  129.6 200.1 132.3 201.3 ;
        RECT  123.3 214.8 134.7 216.0 ;
        RECT  124.5 216.0 125.7 218.1 ;
        RECT  127.5 216.9 128.7 218.1 ;
        RECT  130.5 216.9 131.7 218.1 ;
        RECT  133.5 216.0 134.7 218.1 ;
        RECT  127.2 218.1 128.4 219.0 ;
        RECT  124.5 219.0 125.7 224.7 ;
        RECT  127.2 219.0 129.6 220.2 ;
        RECT  127.2 220.2 128.4 223.5 ;
        RECT  130.8 218.1 132.0 221.7 ;
        RECT  130.2 221.7 132.0 222.9 ;
        RECT  130.8 222.9 132.0 223.5 ;
        RECT  126.9 223.5 128.1 224.7 ;
        RECT  131.1 223.5 132.3 224.7 ;
        RECT  133.5 219.0 134.7 224.7 ;
        RECT  129.0 225.9 130.2 226.2 ;
        RECT  123.3 226.2 134.7 227.4 ;
        RECT  125.4 228.3 128.1 229.5 ;
        RECT  129.6 228.3 132.3 229.5 ;
        RECT  123.3 243.0 134.7 244.2 ;
        RECT  124.5 240.9 125.7 243.0 ;
        RECT  127.5 240.9 128.7 242.1 ;
        RECT  130.5 240.9 131.7 242.1 ;
        RECT  133.5 240.9 134.7 243.0 ;
        RECT  127.2 240.0 128.4 240.9 ;
        RECT  124.5 234.3 125.7 240.0 ;
        RECT  127.2 238.8 129.6 240.0 ;
        RECT  127.2 235.5 128.4 238.8 ;
        RECT  130.8 237.3 132.0 240.9 ;
        RECT  130.2 236.1 132.0 237.3 ;
        RECT  130.8 235.5 132.0 236.1 ;
        RECT  126.9 234.3 128.1 235.5 ;
        RECT  131.1 234.3 132.3 235.5 ;
        RECT  133.5 234.3 134.7 240.0 ;
        RECT  129.0 232.8 130.2 233.1 ;
        RECT  123.3 231.6 134.7 232.8 ;
        RECT  125.4 229.5 128.1 230.7 ;
        RECT  129.6 229.5 132.3 230.7 ;
        RECT  123.3 244.2 134.7 245.4 ;
        RECT  124.5 245.4 125.7 247.5 ;
        RECT  127.5 246.3 128.7 247.5 ;
        RECT  130.5 246.3 131.7 247.5 ;
        RECT  133.5 245.4 134.7 247.5 ;
        RECT  127.2 247.5 128.4 248.4 ;
        RECT  124.5 248.4 125.7 254.1 ;
        RECT  127.2 248.4 129.6 249.6 ;
        RECT  127.2 249.6 128.4 252.9 ;
        RECT  130.8 247.5 132.0 251.1 ;
        RECT  130.2 251.1 132.0 252.3 ;
        RECT  130.8 252.3 132.0 252.9 ;
        RECT  126.9 252.9 128.1 254.1 ;
        RECT  131.1 252.9 132.3 254.1 ;
        RECT  133.5 248.4 134.7 254.1 ;
        RECT  129.0 255.3 130.2 255.6 ;
        RECT  123.3 255.6 134.7 256.8 ;
        RECT  125.4 257.7 128.1 258.9 ;
        RECT  129.6 257.7 132.3 258.9 ;
        RECT  123.3 272.4 134.7 273.6 ;
        RECT  124.5 270.3 125.7 272.4 ;
        RECT  127.5 270.3 128.7 271.5 ;
        RECT  130.5 270.3 131.7 271.5 ;
        RECT  133.5 270.3 134.7 272.4 ;
        RECT  127.2 269.4 128.4 270.3 ;
        RECT  124.5 263.7 125.7 269.4 ;
        RECT  127.2 268.2 129.6 269.4 ;
        RECT  127.2 264.9 128.4 268.2 ;
        RECT  130.8 266.7 132.0 270.3 ;
        RECT  130.2 265.5 132.0 266.7 ;
        RECT  130.8 264.9 132.0 265.5 ;
        RECT  126.9 263.7 128.1 264.9 ;
        RECT  131.1 263.7 132.3 264.9 ;
        RECT  133.5 263.7 134.7 269.4 ;
        RECT  129.0 262.2 130.2 262.5 ;
        RECT  123.3 261.0 134.7 262.2 ;
        RECT  125.4 258.9 128.1 260.1 ;
        RECT  129.6 258.9 132.3 260.1 ;
        RECT  123.3 273.6 134.7 274.8 ;
        RECT  124.5 274.8 125.7 276.9 ;
        RECT  127.5 275.7 128.7 276.9 ;
        RECT  130.5 275.7 131.7 276.9 ;
        RECT  133.5 274.8 134.7 276.9 ;
        RECT  127.2 276.9 128.4 277.8 ;
        RECT  124.5 277.8 125.7 283.5 ;
        RECT  127.2 277.8 129.6 279.0 ;
        RECT  127.2 279.0 128.4 282.3 ;
        RECT  130.8 276.9 132.0 280.5 ;
        RECT  130.2 280.5 132.0 281.7 ;
        RECT  130.8 281.7 132.0 282.3 ;
        RECT  126.9 282.3 128.1 283.5 ;
        RECT  131.1 282.3 132.3 283.5 ;
        RECT  133.5 277.8 134.7 283.5 ;
        RECT  129.0 284.7 130.2 285.0 ;
        RECT  123.3 285.0 134.7 286.2 ;
        RECT  125.4 287.1 128.1 288.3 ;
        RECT  129.6 287.1 132.3 288.3 ;
        RECT  123.3 301.8 134.7 303.0 ;
        RECT  124.5 299.7 125.7 301.8 ;
        RECT  127.5 299.7 128.7 300.9 ;
        RECT  130.5 299.7 131.7 300.9 ;
        RECT  133.5 299.7 134.7 301.8 ;
        RECT  127.2 298.8 128.4 299.7 ;
        RECT  124.5 293.1 125.7 298.8 ;
        RECT  127.2 297.6 129.6 298.8 ;
        RECT  127.2 294.3 128.4 297.6 ;
        RECT  130.8 296.1 132.0 299.7 ;
        RECT  130.2 294.9 132.0 296.1 ;
        RECT  130.8 294.3 132.0 294.9 ;
        RECT  126.9 293.1 128.1 294.3 ;
        RECT  131.1 293.1 132.3 294.3 ;
        RECT  133.5 293.1 134.7 298.8 ;
        RECT  129.0 291.6 130.2 291.9 ;
        RECT  123.3 290.4 134.7 291.6 ;
        RECT  125.4 288.3 128.1 289.5 ;
        RECT  129.6 288.3 132.3 289.5 ;
        RECT  123.3 303.0 134.7 304.2 ;
        RECT  124.5 304.2 125.7 306.3 ;
        RECT  127.5 305.1 128.7 306.3 ;
        RECT  130.5 305.1 131.7 306.3 ;
        RECT  133.5 304.2 134.7 306.3 ;
        RECT  127.2 306.3 128.4 307.2 ;
        RECT  124.5 307.2 125.7 312.9 ;
        RECT  127.2 307.2 129.6 308.4 ;
        RECT  127.2 308.4 128.4 311.7 ;
        RECT  130.8 306.3 132.0 309.9 ;
        RECT  130.2 309.9 132.0 311.1 ;
        RECT  130.8 311.1 132.0 311.7 ;
        RECT  126.9 311.7 128.1 312.9 ;
        RECT  131.1 311.7 132.3 312.9 ;
        RECT  133.5 307.2 134.7 312.9 ;
        RECT  129.0 314.1 130.2 314.4 ;
        RECT  123.3 314.4 134.7 315.6 ;
        RECT  125.4 316.5 128.1 317.7 ;
        RECT  129.6 316.5 132.3 317.7 ;
        RECT  123.3 331.2 134.7 332.4 ;
        RECT  124.5 329.1 125.7 331.2 ;
        RECT  127.5 329.1 128.7 330.3 ;
        RECT  130.5 329.1 131.7 330.3 ;
        RECT  133.5 329.1 134.7 331.2 ;
        RECT  127.2 328.2 128.4 329.1 ;
        RECT  124.5 322.5 125.7 328.2 ;
        RECT  127.2 327.0 129.6 328.2 ;
        RECT  127.2 323.7 128.4 327.0 ;
        RECT  130.8 325.5 132.0 329.1 ;
        RECT  130.2 324.3 132.0 325.5 ;
        RECT  130.8 323.7 132.0 324.3 ;
        RECT  126.9 322.5 128.1 323.7 ;
        RECT  131.1 322.5 132.3 323.7 ;
        RECT  133.5 322.5 134.7 328.2 ;
        RECT  129.0 321.0 130.2 321.3 ;
        RECT  123.3 319.8 134.7 321.0 ;
        RECT  125.4 317.7 128.1 318.9 ;
        RECT  129.6 317.7 132.3 318.9 ;
        RECT  123.3 332.4 134.7 333.6 ;
        RECT  124.5 333.6 125.7 335.7 ;
        RECT  127.5 334.5 128.7 335.7 ;
        RECT  130.5 334.5 131.7 335.7 ;
        RECT  133.5 333.6 134.7 335.7 ;
        RECT  127.2 335.7 128.4 336.6 ;
        RECT  124.5 336.6 125.7 342.3 ;
        RECT  127.2 336.6 129.6 337.8 ;
        RECT  127.2 337.8 128.4 341.1 ;
        RECT  130.8 335.7 132.0 339.3 ;
        RECT  130.2 339.3 132.0 340.5 ;
        RECT  130.8 340.5 132.0 341.1 ;
        RECT  126.9 341.1 128.1 342.3 ;
        RECT  131.1 341.1 132.3 342.3 ;
        RECT  133.5 336.6 134.7 342.3 ;
        RECT  129.0 343.5 130.2 343.8 ;
        RECT  123.3 343.8 134.7 345.0 ;
        RECT  125.4 345.9 128.1 347.1 ;
        RECT  129.6 345.9 132.3 347.1 ;
        RECT  123.3 360.6 134.7 361.8 ;
        RECT  124.5 358.5 125.7 360.6 ;
        RECT  127.5 358.5 128.7 359.7 ;
        RECT  130.5 358.5 131.7 359.7 ;
        RECT  133.5 358.5 134.7 360.6 ;
        RECT  127.2 357.6 128.4 358.5 ;
        RECT  124.5 351.9 125.7 357.6 ;
        RECT  127.2 356.4 129.6 357.6 ;
        RECT  127.2 353.1 128.4 356.4 ;
        RECT  130.8 354.9 132.0 358.5 ;
        RECT  130.2 353.7 132.0 354.9 ;
        RECT  130.8 353.1 132.0 353.7 ;
        RECT  126.9 351.9 128.1 353.1 ;
        RECT  131.1 351.9 132.3 353.1 ;
        RECT  133.5 351.9 134.7 357.6 ;
        RECT  129.0 350.4 130.2 350.7 ;
        RECT  123.3 349.2 134.7 350.4 ;
        RECT  125.4 347.1 128.1 348.3 ;
        RECT  129.6 347.1 132.3 348.3 ;
        RECT  123.3 361.8 134.7 363.0 ;
        RECT  124.5 363.0 125.7 365.1 ;
        RECT  127.5 363.9 128.7 365.1 ;
        RECT  130.5 363.9 131.7 365.1 ;
        RECT  133.5 363.0 134.7 365.1 ;
        RECT  127.2 365.1 128.4 366.0 ;
        RECT  124.5 366.0 125.7 371.7 ;
        RECT  127.2 366.0 129.6 367.2 ;
        RECT  127.2 367.2 128.4 370.5 ;
        RECT  130.8 365.1 132.0 368.7 ;
        RECT  130.2 368.7 132.0 369.9 ;
        RECT  130.8 369.9 132.0 370.5 ;
        RECT  126.9 370.5 128.1 371.7 ;
        RECT  131.1 370.5 132.3 371.7 ;
        RECT  133.5 366.0 134.7 371.7 ;
        RECT  129.0 372.9 130.2 373.2 ;
        RECT  123.3 373.2 134.7 374.4 ;
        RECT  125.4 375.3 128.1 376.5 ;
        RECT  129.6 375.3 132.3 376.5 ;
        RECT  123.3 390.0 134.7 391.2 ;
        RECT  124.5 387.9 125.7 390.0 ;
        RECT  127.5 387.9 128.7 389.1 ;
        RECT  130.5 387.9 131.7 389.1 ;
        RECT  133.5 387.9 134.7 390.0 ;
        RECT  127.2 387.0 128.4 387.9 ;
        RECT  124.5 381.3 125.7 387.0 ;
        RECT  127.2 385.8 129.6 387.0 ;
        RECT  127.2 382.5 128.4 385.8 ;
        RECT  130.8 384.3 132.0 387.9 ;
        RECT  130.2 383.1 132.0 384.3 ;
        RECT  130.8 382.5 132.0 383.1 ;
        RECT  126.9 381.3 128.1 382.5 ;
        RECT  131.1 381.3 132.3 382.5 ;
        RECT  133.5 381.3 134.7 387.0 ;
        RECT  129.0 379.8 130.2 380.1 ;
        RECT  123.3 378.6 134.7 379.8 ;
        RECT  125.4 376.5 128.1 377.7 ;
        RECT  129.6 376.5 132.3 377.7 ;
        RECT  123.3 391.2 134.7 392.4 ;
        RECT  124.5 392.4 125.7 394.5 ;
        RECT  127.5 393.3 128.7 394.5 ;
        RECT  130.5 393.3 131.7 394.5 ;
        RECT  133.5 392.4 134.7 394.5 ;
        RECT  127.2 394.5 128.4 395.4 ;
        RECT  124.5 395.4 125.7 401.1 ;
        RECT  127.2 395.4 129.6 396.6 ;
        RECT  127.2 396.6 128.4 399.9 ;
        RECT  130.8 394.5 132.0 398.1 ;
        RECT  130.2 398.1 132.0 399.3 ;
        RECT  130.8 399.3 132.0 399.9 ;
        RECT  126.9 399.9 128.1 401.1 ;
        RECT  131.1 399.9 132.3 401.1 ;
        RECT  133.5 395.4 134.7 401.1 ;
        RECT  129.0 402.3 130.2 402.6 ;
        RECT  123.3 402.6 134.7 403.8 ;
        RECT  125.4 404.7 128.1 405.9 ;
        RECT  129.6 404.7 132.3 405.9 ;
        RECT  123.3 419.4 134.7 420.6 ;
        RECT  124.5 417.3 125.7 419.4 ;
        RECT  127.5 417.3 128.7 418.5 ;
        RECT  130.5 417.3 131.7 418.5 ;
        RECT  133.5 417.3 134.7 419.4 ;
        RECT  127.2 416.4 128.4 417.3 ;
        RECT  124.5 410.7 125.7 416.4 ;
        RECT  127.2 415.2 129.6 416.4 ;
        RECT  127.2 411.9 128.4 415.2 ;
        RECT  130.8 413.7 132.0 417.3 ;
        RECT  130.2 412.5 132.0 413.7 ;
        RECT  130.8 411.9 132.0 412.5 ;
        RECT  126.9 410.7 128.1 411.9 ;
        RECT  131.1 410.7 132.3 411.9 ;
        RECT  133.5 410.7 134.7 416.4 ;
        RECT  129.0 409.2 130.2 409.5 ;
        RECT  123.3 408.0 134.7 409.2 ;
        RECT  125.4 405.9 128.1 407.1 ;
        RECT  129.6 405.9 132.3 407.1 ;
        RECT  123.3 420.6 134.7 421.8 ;
        RECT  124.5 421.8 125.7 423.9 ;
        RECT  127.5 422.7 128.7 423.9 ;
        RECT  130.5 422.7 131.7 423.9 ;
        RECT  133.5 421.8 134.7 423.9 ;
        RECT  127.2 423.9 128.4 424.8 ;
        RECT  124.5 424.8 125.7 430.5 ;
        RECT  127.2 424.8 129.6 426.0 ;
        RECT  127.2 426.0 128.4 429.3 ;
        RECT  130.8 423.9 132.0 427.5 ;
        RECT  130.2 427.5 132.0 428.7 ;
        RECT  130.8 428.7 132.0 429.3 ;
        RECT  126.9 429.3 128.1 430.5 ;
        RECT  131.1 429.3 132.3 430.5 ;
        RECT  133.5 424.8 134.7 430.5 ;
        RECT  129.0 431.7 130.2 432.0 ;
        RECT  123.3 432.0 134.7 433.2 ;
        RECT  125.4 434.1 128.1 435.3 ;
        RECT  129.6 434.1 132.3 435.3 ;
        RECT  133.5 213.6 144.9 214.8 ;
        RECT  134.7 211.5 135.9 213.6 ;
        RECT  137.7 211.5 138.9 212.7 ;
        RECT  140.7 211.5 141.9 212.7 ;
        RECT  143.7 211.5 144.9 213.6 ;
        RECT  137.4 210.6 138.6 211.5 ;
        RECT  134.7 204.9 135.9 210.6 ;
        RECT  137.4 209.4 139.8 210.6 ;
        RECT  137.4 206.1 138.6 209.4 ;
        RECT  141.0 207.9 142.2 211.5 ;
        RECT  140.4 206.7 142.2 207.9 ;
        RECT  141.0 206.1 142.2 206.7 ;
        RECT  137.1 204.9 138.3 206.1 ;
        RECT  141.3 204.9 142.5 206.1 ;
        RECT  143.7 204.9 144.9 210.6 ;
        RECT  139.2 203.4 140.4 203.7 ;
        RECT  133.5 202.2 144.9 203.4 ;
        RECT  135.6 200.1 138.3 201.3 ;
        RECT  139.8 200.1 142.5 201.3 ;
        RECT  133.5 214.8 144.9 216.0 ;
        RECT  134.7 216.0 135.9 218.1 ;
        RECT  137.7 216.9 138.9 218.1 ;
        RECT  140.7 216.9 141.9 218.1 ;
        RECT  143.7 216.0 144.9 218.1 ;
        RECT  137.4 218.1 138.6 219.0 ;
        RECT  134.7 219.0 135.9 224.7 ;
        RECT  137.4 219.0 139.8 220.2 ;
        RECT  137.4 220.2 138.6 223.5 ;
        RECT  141.0 218.1 142.2 221.7 ;
        RECT  140.4 221.7 142.2 222.9 ;
        RECT  141.0 222.9 142.2 223.5 ;
        RECT  137.1 223.5 138.3 224.7 ;
        RECT  141.3 223.5 142.5 224.7 ;
        RECT  143.7 219.0 144.9 224.7 ;
        RECT  139.2 225.9 140.4 226.2 ;
        RECT  133.5 226.2 144.9 227.4 ;
        RECT  135.6 228.3 138.3 229.5 ;
        RECT  139.8 228.3 142.5 229.5 ;
        RECT  133.5 243.0 144.9 244.2 ;
        RECT  134.7 240.9 135.9 243.0 ;
        RECT  137.7 240.9 138.9 242.1 ;
        RECT  140.7 240.9 141.9 242.1 ;
        RECT  143.7 240.9 144.9 243.0 ;
        RECT  137.4 240.0 138.6 240.9 ;
        RECT  134.7 234.3 135.9 240.0 ;
        RECT  137.4 238.8 139.8 240.0 ;
        RECT  137.4 235.5 138.6 238.8 ;
        RECT  141.0 237.3 142.2 240.9 ;
        RECT  140.4 236.1 142.2 237.3 ;
        RECT  141.0 235.5 142.2 236.1 ;
        RECT  137.1 234.3 138.3 235.5 ;
        RECT  141.3 234.3 142.5 235.5 ;
        RECT  143.7 234.3 144.9 240.0 ;
        RECT  139.2 232.8 140.4 233.1 ;
        RECT  133.5 231.6 144.9 232.8 ;
        RECT  135.6 229.5 138.3 230.7 ;
        RECT  139.8 229.5 142.5 230.7 ;
        RECT  133.5 244.2 144.9 245.4 ;
        RECT  134.7 245.4 135.9 247.5 ;
        RECT  137.7 246.3 138.9 247.5 ;
        RECT  140.7 246.3 141.9 247.5 ;
        RECT  143.7 245.4 144.9 247.5 ;
        RECT  137.4 247.5 138.6 248.4 ;
        RECT  134.7 248.4 135.9 254.1 ;
        RECT  137.4 248.4 139.8 249.6 ;
        RECT  137.4 249.6 138.6 252.9 ;
        RECT  141.0 247.5 142.2 251.1 ;
        RECT  140.4 251.1 142.2 252.3 ;
        RECT  141.0 252.3 142.2 252.9 ;
        RECT  137.1 252.9 138.3 254.1 ;
        RECT  141.3 252.9 142.5 254.1 ;
        RECT  143.7 248.4 144.9 254.1 ;
        RECT  139.2 255.3 140.4 255.6 ;
        RECT  133.5 255.6 144.9 256.8 ;
        RECT  135.6 257.7 138.3 258.9 ;
        RECT  139.8 257.7 142.5 258.9 ;
        RECT  133.5 272.4 144.9 273.6 ;
        RECT  134.7 270.3 135.9 272.4 ;
        RECT  137.7 270.3 138.9 271.5 ;
        RECT  140.7 270.3 141.9 271.5 ;
        RECT  143.7 270.3 144.9 272.4 ;
        RECT  137.4 269.4 138.6 270.3 ;
        RECT  134.7 263.7 135.9 269.4 ;
        RECT  137.4 268.2 139.8 269.4 ;
        RECT  137.4 264.9 138.6 268.2 ;
        RECT  141.0 266.7 142.2 270.3 ;
        RECT  140.4 265.5 142.2 266.7 ;
        RECT  141.0 264.9 142.2 265.5 ;
        RECT  137.1 263.7 138.3 264.9 ;
        RECT  141.3 263.7 142.5 264.9 ;
        RECT  143.7 263.7 144.9 269.4 ;
        RECT  139.2 262.2 140.4 262.5 ;
        RECT  133.5 261.0 144.9 262.2 ;
        RECT  135.6 258.9 138.3 260.1 ;
        RECT  139.8 258.9 142.5 260.1 ;
        RECT  133.5 273.6 144.9 274.8 ;
        RECT  134.7 274.8 135.9 276.9 ;
        RECT  137.7 275.7 138.9 276.9 ;
        RECT  140.7 275.7 141.9 276.9 ;
        RECT  143.7 274.8 144.9 276.9 ;
        RECT  137.4 276.9 138.6 277.8 ;
        RECT  134.7 277.8 135.9 283.5 ;
        RECT  137.4 277.8 139.8 279.0 ;
        RECT  137.4 279.0 138.6 282.3 ;
        RECT  141.0 276.9 142.2 280.5 ;
        RECT  140.4 280.5 142.2 281.7 ;
        RECT  141.0 281.7 142.2 282.3 ;
        RECT  137.1 282.3 138.3 283.5 ;
        RECT  141.3 282.3 142.5 283.5 ;
        RECT  143.7 277.8 144.9 283.5 ;
        RECT  139.2 284.7 140.4 285.0 ;
        RECT  133.5 285.0 144.9 286.2 ;
        RECT  135.6 287.1 138.3 288.3 ;
        RECT  139.8 287.1 142.5 288.3 ;
        RECT  133.5 301.8 144.9 303.0 ;
        RECT  134.7 299.7 135.9 301.8 ;
        RECT  137.7 299.7 138.9 300.9 ;
        RECT  140.7 299.7 141.9 300.9 ;
        RECT  143.7 299.7 144.9 301.8 ;
        RECT  137.4 298.8 138.6 299.7 ;
        RECT  134.7 293.1 135.9 298.8 ;
        RECT  137.4 297.6 139.8 298.8 ;
        RECT  137.4 294.3 138.6 297.6 ;
        RECT  141.0 296.1 142.2 299.7 ;
        RECT  140.4 294.9 142.2 296.1 ;
        RECT  141.0 294.3 142.2 294.9 ;
        RECT  137.1 293.1 138.3 294.3 ;
        RECT  141.3 293.1 142.5 294.3 ;
        RECT  143.7 293.1 144.9 298.8 ;
        RECT  139.2 291.6 140.4 291.9 ;
        RECT  133.5 290.4 144.9 291.6 ;
        RECT  135.6 288.3 138.3 289.5 ;
        RECT  139.8 288.3 142.5 289.5 ;
        RECT  133.5 303.0 144.9 304.2 ;
        RECT  134.7 304.2 135.9 306.3 ;
        RECT  137.7 305.1 138.9 306.3 ;
        RECT  140.7 305.1 141.9 306.3 ;
        RECT  143.7 304.2 144.9 306.3 ;
        RECT  137.4 306.3 138.6 307.2 ;
        RECT  134.7 307.2 135.9 312.9 ;
        RECT  137.4 307.2 139.8 308.4 ;
        RECT  137.4 308.4 138.6 311.7 ;
        RECT  141.0 306.3 142.2 309.9 ;
        RECT  140.4 309.9 142.2 311.1 ;
        RECT  141.0 311.1 142.2 311.7 ;
        RECT  137.1 311.7 138.3 312.9 ;
        RECT  141.3 311.7 142.5 312.9 ;
        RECT  143.7 307.2 144.9 312.9 ;
        RECT  139.2 314.1 140.4 314.4 ;
        RECT  133.5 314.4 144.9 315.6 ;
        RECT  135.6 316.5 138.3 317.7 ;
        RECT  139.8 316.5 142.5 317.7 ;
        RECT  133.5 331.2 144.9 332.4 ;
        RECT  134.7 329.1 135.9 331.2 ;
        RECT  137.7 329.1 138.9 330.3 ;
        RECT  140.7 329.1 141.9 330.3 ;
        RECT  143.7 329.1 144.9 331.2 ;
        RECT  137.4 328.2 138.6 329.1 ;
        RECT  134.7 322.5 135.9 328.2 ;
        RECT  137.4 327.0 139.8 328.2 ;
        RECT  137.4 323.7 138.6 327.0 ;
        RECT  141.0 325.5 142.2 329.1 ;
        RECT  140.4 324.3 142.2 325.5 ;
        RECT  141.0 323.7 142.2 324.3 ;
        RECT  137.1 322.5 138.3 323.7 ;
        RECT  141.3 322.5 142.5 323.7 ;
        RECT  143.7 322.5 144.9 328.2 ;
        RECT  139.2 321.0 140.4 321.3 ;
        RECT  133.5 319.8 144.9 321.0 ;
        RECT  135.6 317.7 138.3 318.9 ;
        RECT  139.8 317.7 142.5 318.9 ;
        RECT  133.5 332.4 144.9 333.6 ;
        RECT  134.7 333.6 135.9 335.7 ;
        RECT  137.7 334.5 138.9 335.7 ;
        RECT  140.7 334.5 141.9 335.7 ;
        RECT  143.7 333.6 144.9 335.7 ;
        RECT  137.4 335.7 138.6 336.6 ;
        RECT  134.7 336.6 135.9 342.3 ;
        RECT  137.4 336.6 139.8 337.8 ;
        RECT  137.4 337.8 138.6 341.1 ;
        RECT  141.0 335.7 142.2 339.3 ;
        RECT  140.4 339.3 142.2 340.5 ;
        RECT  141.0 340.5 142.2 341.1 ;
        RECT  137.1 341.1 138.3 342.3 ;
        RECT  141.3 341.1 142.5 342.3 ;
        RECT  143.7 336.6 144.9 342.3 ;
        RECT  139.2 343.5 140.4 343.8 ;
        RECT  133.5 343.8 144.9 345.0 ;
        RECT  135.6 345.9 138.3 347.1 ;
        RECT  139.8 345.9 142.5 347.1 ;
        RECT  133.5 360.6 144.9 361.8 ;
        RECT  134.7 358.5 135.9 360.6 ;
        RECT  137.7 358.5 138.9 359.7 ;
        RECT  140.7 358.5 141.9 359.7 ;
        RECT  143.7 358.5 144.9 360.6 ;
        RECT  137.4 357.6 138.6 358.5 ;
        RECT  134.7 351.9 135.9 357.6 ;
        RECT  137.4 356.4 139.8 357.6 ;
        RECT  137.4 353.1 138.6 356.4 ;
        RECT  141.0 354.9 142.2 358.5 ;
        RECT  140.4 353.7 142.2 354.9 ;
        RECT  141.0 353.1 142.2 353.7 ;
        RECT  137.1 351.9 138.3 353.1 ;
        RECT  141.3 351.9 142.5 353.1 ;
        RECT  143.7 351.9 144.9 357.6 ;
        RECT  139.2 350.4 140.4 350.7 ;
        RECT  133.5 349.2 144.9 350.4 ;
        RECT  135.6 347.1 138.3 348.3 ;
        RECT  139.8 347.1 142.5 348.3 ;
        RECT  133.5 361.8 144.9 363.0 ;
        RECT  134.7 363.0 135.9 365.1 ;
        RECT  137.7 363.9 138.9 365.1 ;
        RECT  140.7 363.9 141.9 365.1 ;
        RECT  143.7 363.0 144.9 365.1 ;
        RECT  137.4 365.1 138.6 366.0 ;
        RECT  134.7 366.0 135.9 371.7 ;
        RECT  137.4 366.0 139.8 367.2 ;
        RECT  137.4 367.2 138.6 370.5 ;
        RECT  141.0 365.1 142.2 368.7 ;
        RECT  140.4 368.7 142.2 369.9 ;
        RECT  141.0 369.9 142.2 370.5 ;
        RECT  137.1 370.5 138.3 371.7 ;
        RECT  141.3 370.5 142.5 371.7 ;
        RECT  143.7 366.0 144.9 371.7 ;
        RECT  139.2 372.9 140.4 373.2 ;
        RECT  133.5 373.2 144.9 374.4 ;
        RECT  135.6 375.3 138.3 376.5 ;
        RECT  139.8 375.3 142.5 376.5 ;
        RECT  133.5 390.0 144.9 391.2 ;
        RECT  134.7 387.9 135.9 390.0 ;
        RECT  137.7 387.9 138.9 389.1 ;
        RECT  140.7 387.9 141.9 389.1 ;
        RECT  143.7 387.9 144.9 390.0 ;
        RECT  137.4 387.0 138.6 387.9 ;
        RECT  134.7 381.3 135.9 387.0 ;
        RECT  137.4 385.8 139.8 387.0 ;
        RECT  137.4 382.5 138.6 385.8 ;
        RECT  141.0 384.3 142.2 387.9 ;
        RECT  140.4 383.1 142.2 384.3 ;
        RECT  141.0 382.5 142.2 383.1 ;
        RECT  137.1 381.3 138.3 382.5 ;
        RECT  141.3 381.3 142.5 382.5 ;
        RECT  143.7 381.3 144.9 387.0 ;
        RECT  139.2 379.8 140.4 380.1 ;
        RECT  133.5 378.6 144.9 379.8 ;
        RECT  135.6 376.5 138.3 377.7 ;
        RECT  139.8 376.5 142.5 377.7 ;
        RECT  133.5 391.2 144.9 392.4 ;
        RECT  134.7 392.4 135.9 394.5 ;
        RECT  137.7 393.3 138.9 394.5 ;
        RECT  140.7 393.3 141.9 394.5 ;
        RECT  143.7 392.4 144.9 394.5 ;
        RECT  137.4 394.5 138.6 395.4 ;
        RECT  134.7 395.4 135.9 401.1 ;
        RECT  137.4 395.4 139.8 396.6 ;
        RECT  137.4 396.6 138.6 399.9 ;
        RECT  141.0 394.5 142.2 398.1 ;
        RECT  140.4 398.1 142.2 399.3 ;
        RECT  141.0 399.3 142.2 399.9 ;
        RECT  137.1 399.9 138.3 401.1 ;
        RECT  141.3 399.9 142.5 401.1 ;
        RECT  143.7 395.4 144.9 401.1 ;
        RECT  139.2 402.3 140.4 402.6 ;
        RECT  133.5 402.6 144.9 403.8 ;
        RECT  135.6 404.7 138.3 405.9 ;
        RECT  139.8 404.7 142.5 405.9 ;
        RECT  133.5 419.4 144.9 420.6 ;
        RECT  134.7 417.3 135.9 419.4 ;
        RECT  137.7 417.3 138.9 418.5 ;
        RECT  140.7 417.3 141.9 418.5 ;
        RECT  143.7 417.3 144.9 419.4 ;
        RECT  137.4 416.4 138.6 417.3 ;
        RECT  134.7 410.7 135.9 416.4 ;
        RECT  137.4 415.2 139.8 416.4 ;
        RECT  137.4 411.9 138.6 415.2 ;
        RECT  141.0 413.7 142.2 417.3 ;
        RECT  140.4 412.5 142.2 413.7 ;
        RECT  141.0 411.9 142.2 412.5 ;
        RECT  137.1 410.7 138.3 411.9 ;
        RECT  141.3 410.7 142.5 411.9 ;
        RECT  143.7 410.7 144.9 416.4 ;
        RECT  139.2 409.2 140.4 409.5 ;
        RECT  133.5 408.0 144.9 409.2 ;
        RECT  135.6 405.9 138.3 407.1 ;
        RECT  139.8 405.9 142.5 407.1 ;
        RECT  133.5 420.6 144.9 421.8 ;
        RECT  134.7 421.8 135.9 423.9 ;
        RECT  137.7 422.7 138.9 423.9 ;
        RECT  140.7 422.7 141.9 423.9 ;
        RECT  143.7 421.8 144.9 423.9 ;
        RECT  137.4 423.9 138.6 424.8 ;
        RECT  134.7 424.8 135.9 430.5 ;
        RECT  137.4 424.8 139.8 426.0 ;
        RECT  137.4 426.0 138.6 429.3 ;
        RECT  141.0 423.9 142.2 427.5 ;
        RECT  140.4 427.5 142.2 428.7 ;
        RECT  141.0 428.7 142.2 429.3 ;
        RECT  137.1 429.3 138.3 430.5 ;
        RECT  141.3 429.3 142.5 430.5 ;
        RECT  143.7 424.8 144.9 430.5 ;
        RECT  139.2 431.7 140.4 432.0 ;
        RECT  133.5 432.0 144.9 433.2 ;
        RECT  135.6 434.1 138.3 435.3 ;
        RECT  139.8 434.1 142.5 435.3 ;
        RECT  143.7 213.6 155.1 214.8 ;
        RECT  144.9 211.5 146.1 213.6 ;
        RECT  147.9 211.5 149.1 212.7 ;
        RECT  150.9 211.5 152.1 212.7 ;
        RECT  153.9 211.5 155.1 213.6 ;
        RECT  147.6 210.6 148.8 211.5 ;
        RECT  144.9 204.9 146.1 210.6 ;
        RECT  147.6 209.4 150.0 210.6 ;
        RECT  147.6 206.1 148.8 209.4 ;
        RECT  151.2 207.9 152.4 211.5 ;
        RECT  150.6 206.7 152.4 207.9 ;
        RECT  151.2 206.1 152.4 206.7 ;
        RECT  147.3 204.9 148.5 206.1 ;
        RECT  151.5 204.9 152.7 206.1 ;
        RECT  153.9 204.9 155.1 210.6 ;
        RECT  149.4 203.4 150.6 203.7 ;
        RECT  143.7 202.2 155.1 203.4 ;
        RECT  145.8 200.1 148.5 201.3 ;
        RECT  150.0 200.1 152.7 201.3 ;
        RECT  143.7 214.8 155.1 216.0 ;
        RECT  144.9 216.0 146.1 218.1 ;
        RECT  147.9 216.9 149.1 218.1 ;
        RECT  150.9 216.9 152.1 218.1 ;
        RECT  153.9 216.0 155.1 218.1 ;
        RECT  147.6 218.1 148.8 219.0 ;
        RECT  144.9 219.0 146.1 224.7 ;
        RECT  147.6 219.0 150.0 220.2 ;
        RECT  147.6 220.2 148.8 223.5 ;
        RECT  151.2 218.1 152.4 221.7 ;
        RECT  150.6 221.7 152.4 222.9 ;
        RECT  151.2 222.9 152.4 223.5 ;
        RECT  147.3 223.5 148.5 224.7 ;
        RECT  151.5 223.5 152.7 224.7 ;
        RECT  153.9 219.0 155.1 224.7 ;
        RECT  149.4 225.9 150.6 226.2 ;
        RECT  143.7 226.2 155.1 227.4 ;
        RECT  145.8 228.3 148.5 229.5 ;
        RECT  150.0 228.3 152.7 229.5 ;
        RECT  143.7 243.0 155.1 244.2 ;
        RECT  144.9 240.9 146.1 243.0 ;
        RECT  147.9 240.9 149.1 242.1 ;
        RECT  150.9 240.9 152.1 242.1 ;
        RECT  153.9 240.9 155.1 243.0 ;
        RECT  147.6 240.0 148.8 240.9 ;
        RECT  144.9 234.3 146.1 240.0 ;
        RECT  147.6 238.8 150.0 240.0 ;
        RECT  147.6 235.5 148.8 238.8 ;
        RECT  151.2 237.3 152.4 240.9 ;
        RECT  150.6 236.1 152.4 237.3 ;
        RECT  151.2 235.5 152.4 236.1 ;
        RECT  147.3 234.3 148.5 235.5 ;
        RECT  151.5 234.3 152.7 235.5 ;
        RECT  153.9 234.3 155.1 240.0 ;
        RECT  149.4 232.8 150.6 233.1 ;
        RECT  143.7 231.6 155.1 232.8 ;
        RECT  145.8 229.5 148.5 230.7 ;
        RECT  150.0 229.5 152.7 230.7 ;
        RECT  143.7 244.2 155.1 245.4 ;
        RECT  144.9 245.4 146.1 247.5 ;
        RECT  147.9 246.3 149.1 247.5 ;
        RECT  150.9 246.3 152.1 247.5 ;
        RECT  153.9 245.4 155.1 247.5 ;
        RECT  147.6 247.5 148.8 248.4 ;
        RECT  144.9 248.4 146.1 254.1 ;
        RECT  147.6 248.4 150.0 249.6 ;
        RECT  147.6 249.6 148.8 252.9 ;
        RECT  151.2 247.5 152.4 251.1 ;
        RECT  150.6 251.1 152.4 252.3 ;
        RECT  151.2 252.3 152.4 252.9 ;
        RECT  147.3 252.9 148.5 254.1 ;
        RECT  151.5 252.9 152.7 254.1 ;
        RECT  153.9 248.4 155.1 254.1 ;
        RECT  149.4 255.3 150.6 255.6 ;
        RECT  143.7 255.6 155.1 256.8 ;
        RECT  145.8 257.7 148.5 258.9 ;
        RECT  150.0 257.7 152.7 258.9 ;
        RECT  143.7 272.4 155.1 273.6 ;
        RECT  144.9 270.3 146.1 272.4 ;
        RECT  147.9 270.3 149.1 271.5 ;
        RECT  150.9 270.3 152.1 271.5 ;
        RECT  153.9 270.3 155.1 272.4 ;
        RECT  147.6 269.4 148.8 270.3 ;
        RECT  144.9 263.7 146.1 269.4 ;
        RECT  147.6 268.2 150.0 269.4 ;
        RECT  147.6 264.9 148.8 268.2 ;
        RECT  151.2 266.7 152.4 270.3 ;
        RECT  150.6 265.5 152.4 266.7 ;
        RECT  151.2 264.9 152.4 265.5 ;
        RECT  147.3 263.7 148.5 264.9 ;
        RECT  151.5 263.7 152.7 264.9 ;
        RECT  153.9 263.7 155.1 269.4 ;
        RECT  149.4 262.2 150.6 262.5 ;
        RECT  143.7 261.0 155.1 262.2 ;
        RECT  145.8 258.9 148.5 260.1 ;
        RECT  150.0 258.9 152.7 260.1 ;
        RECT  143.7 273.6 155.1 274.8 ;
        RECT  144.9 274.8 146.1 276.9 ;
        RECT  147.9 275.7 149.1 276.9 ;
        RECT  150.9 275.7 152.1 276.9 ;
        RECT  153.9 274.8 155.1 276.9 ;
        RECT  147.6 276.9 148.8 277.8 ;
        RECT  144.9 277.8 146.1 283.5 ;
        RECT  147.6 277.8 150.0 279.0 ;
        RECT  147.6 279.0 148.8 282.3 ;
        RECT  151.2 276.9 152.4 280.5 ;
        RECT  150.6 280.5 152.4 281.7 ;
        RECT  151.2 281.7 152.4 282.3 ;
        RECT  147.3 282.3 148.5 283.5 ;
        RECT  151.5 282.3 152.7 283.5 ;
        RECT  153.9 277.8 155.1 283.5 ;
        RECT  149.4 284.7 150.6 285.0 ;
        RECT  143.7 285.0 155.1 286.2 ;
        RECT  145.8 287.1 148.5 288.3 ;
        RECT  150.0 287.1 152.7 288.3 ;
        RECT  143.7 301.8 155.1 303.0 ;
        RECT  144.9 299.7 146.1 301.8 ;
        RECT  147.9 299.7 149.1 300.9 ;
        RECT  150.9 299.7 152.1 300.9 ;
        RECT  153.9 299.7 155.1 301.8 ;
        RECT  147.6 298.8 148.8 299.7 ;
        RECT  144.9 293.1 146.1 298.8 ;
        RECT  147.6 297.6 150.0 298.8 ;
        RECT  147.6 294.3 148.8 297.6 ;
        RECT  151.2 296.1 152.4 299.7 ;
        RECT  150.6 294.9 152.4 296.1 ;
        RECT  151.2 294.3 152.4 294.9 ;
        RECT  147.3 293.1 148.5 294.3 ;
        RECT  151.5 293.1 152.7 294.3 ;
        RECT  153.9 293.1 155.1 298.8 ;
        RECT  149.4 291.6 150.6 291.9 ;
        RECT  143.7 290.4 155.1 291.6 ;
        RECT  145.8 288.3 148.5 289.5 ;
        RECT  150.0 288.3 152.7 289.5 ;
        RECT  143.7 303.0 155.1 304.2 ;
        RECT  144.9 304.2 146.1 306.3 ;
        RECT  147.9 305.1 149.1 306.3 ;
        RECT  150.9 305.1 152.1 306.3 ;
        RECT  153.9 304.2 155.1 306.3 ;
        RECT  147.6 306.3 148.8 307.2 ;
        RECT  144.9 307.2 146.1 312.9 ;
        RECT  147.6 307.2 150.0 308.4 ;
        RECT  147.6 308.4 148.8 311.7 ;
        RECT  151.2 306.3 152.4 309.9 ;
        RECT  150.6 309.9 152.4 311.1 ;
        RECT  151.2 311.1 152.4 311.7 ;
        RECT  147.3 311.7 148.5 312.9 ;
        RECT  151.5 311.7 152.7 312.9 ;
        RECT  153.9 307.2 155.1 312.9 ;
        RECT  149.4 314.1 150.6 314.4 ;
        RECT  143.7 314.4 155.1 315.6 ;
        RECT  145.8 316.5 148.5 317.7 ;
        RECT  150.0 316.5 152.7 317.7 ;
        RECT  143.7 331.2 155.1 332.4 ;
        RECT  144.9 329.1 146.1 331.2 ;
        RECT  147.9 329.1 149.1 330.3 ;
        RECT  150.9 329.1 152.1 330.3 ;
        RECT  153.9 329.1 155.1 331.2 ;
        RECT  147.6 328.2 148.8 329.1 ;
        RECT  144.9 322.5 146.1 328.2 ;
        RECT  147.6 327.0 150.0 328.2 ;
        RECT  147.6 323.7 148.8 327.0 ;
        RECT  151.2 325.5 152.4 329.1 ;
        RECT  150.6 324.3 152.4 325.5 ;
        RECT  151.2 323.7 152.4 324.3 ;
        RECT  147.3 322.5 148.5 323.7 ;
        RECT  151.5 322.5 152.7 323.7 ;
        RECT  153.9 322.5 155.1 328.2 ;
        RECT  149.4 321.0 150.6 321.3 ;
        RECT  143.7 319.8 155.1 321.0 ;
        RECT  145.8 317.7 148.5 318.9 ;
        RECT  150.0 317.7 152.7 318.9 ;
        RECT  143.7 332.4 155.1 333.6 ;
        RECT  144.9 333.6 146.1 335.7 ;
        RECT  147.9 334.5 149.1 335.7 ;
        RECT  150.9 334.5 152.1 335.7 ;
        RECT  153.9 333.6 155.1 335.7 ;
        RECT  147.6 335.7 148.8 336.6 ;
        RECT  144.9 336.6 146.1 342.3 ;
        RECT  147.6 336.6 150.0 337.8 ;
        RECT  147.6 337.8 148.8 341.1 ;
        RECT  151.2 335.7 152.4 339.3 ;
        RECT  150.6 339.3 152.4 340.5 ;
        RECT  151.2 340.5 152.4 341.1 ;
        RECT  147.3 341.1 148.5 342.3 ;
        RECT  151.5 341.1 152.7 342.3 ;
        RECT  153.9 336.6 155.1 342.3 ;
        RECT  149.4 343.5 150.6 343.8 ;
        RECT  143.7 343.8 155.1 345.0 ;
        RECT  145.8 345.9 148.5 347.1 ;
        RECT  150.0 345.9 152.7 347.1 ;
        RECT  143.7 360.6 155.1 361.8 ;
        RECT  144.9 358.5 146.1 360.6 ;
        RECT  147.9 358.5 149.1 359.7 ;
        RECT  150.9 358.5 152.1 359.7 ;
        RECT  153.9 358.5 155.1 360.6 ;
        RECT  147.6 357.6 148.8 358.5 ;
        RECT  144.9 351.9 146.1 357.6 ;
        RECT  147.6 356.4 150.0 357.6 ;
        RECT  147.6 353.1 148.8 356.4 ;
        RECT  151.2 354.9 152.4 358.5 ;
        RECT  150.6 353.7 152.4 354.9 ;
        RECT  151.2 353.1 152.4 353.7 ;
        RECT  147.3 351.9 148.5 353.1 ;
        RECT  151.5 351.9 152.7 353.1 ;
        RECT  153.9 351.9 155.1 357.6 ;
        RECT  149.4 350.4 150.6 350.7 ;
        RECT  143.7 349.2 155.1 350.4 ;
        RECT  145.8 347.1 148.5 348.3 ;
        RECT  150.0 347.1 152.7 348.3 ;
        RECT  143.7 361.8 155.1 363.0 ;
        RECT  144.9 363.0 146.1 365.1 ;
        RECT  147.9 363.9 149.1 365.1 ;
        RECT  150.9 363.9 152.1 365.1 ;
        RECT  153.9 363.0 155.1 365.1 ;
        RECT  147.6 365.1 148.8 366.0 ;
        RECT  144.9 366.0 146.1 371.7 ;
        RECT  147.6 366.0 150.0 367.2 ;
        RECT  147.6 367.2 148.8 370.5 ;
        RECT  151.2 365.1 152.4 368.7 ;
        RECT  150.6 368.7 152.4 369.9 ;
        RECT  151.2 369.9 152.4 370.5 ;
        RECT  147.3 370.5 148.5 371.7 ;
        RECT  151.5 370.5 152.7 371.7 ;
        RECT  153.9 366.0 155.1 371.7 ;
        RECT  149.4 372.9 150.6 373.2 ;
        RECT  143.7 373.2 155.1 374.4 ;
        RECT  145.8 375.3 148.5 376.5 ;
        RECT  150.0 375.3 152.7 376.5 ;
        RECT  143.7 390.0 155.1 391.2 ;
        RECT  144.9 387.9 146.1 390.0 ;
        RECT  147.9 387.9 149.1 389.1 ;
        RECT  150.9 387.9 152.1 389.1 ;
        RECT  153.9 387.9 155.1 390.0 ;
        RECT  147.6 387.0 148.8 387.9 ;
        RECT  144.9 381.3 146.1 387.0 ;
        RECT  147.6 385.8 150.0 387.0 ;
        RECT  147.6 382.5 148.8 385.8 ;
        RECT  151.2 384.3 152.4 387.9 ;
        RECT  150.6 383.1 152.4 384.3 ;
        RECT  151.2 382.5 152.4 383.1 ;
        RECT  147.3 381.3 148.5 382.5 ;
        RECT  151.5 381.3 152.7 382.5 ;
        RECT  153.9 381.3 155.1 387.0 ;
        RECT  149.4 379.8 150.6 380.1 ;
        RECT  143.7 378.6 155.1 379.8 ;
        RECT  145.8 376.5 148.5 377.7 ;
        RECT  150.0 376.5 152.7 377.7 ;
        RECT  143.7 391.2 155.1 392.4 ;
        RECT  144.9 392.4 146.1 394.5 ;
        RECT  147.9 393.3 149.1 394.5 ;
        RECT  150.9 393.3 152.1 394.5 ;
        RECT  153.9 392.4 155.1 394.5 ;
        RECT  147.6 394.5 148.8 395.4 ;
        RECT  144.9 395.4 146.1 401.1 ;
        RECT  147.6 395.4 150.0 396.6 ;
        RECT  147.6 396.6 148.8 399.9 ;
        RECT  151.2 394.5 152.4 398.1 ;
        RECT  150.6 398.1 152.4 399.3 ;
        RECT  151.2 399.3 152.4 399.9 ;
        RECT  147.3 399.9 148.5 401.1 ;
        RECT  151.5 399.9 152.7 401.1 ;
        RECT  153.9 395.4 155.1 401.1 ;
        RECT  149.4 402.3 150.6 402.6 ;
        RECT  143.7 402.6 155.1 403.8 ;
        RECT  145.8 404.7 148.5 405.9 ;
        RECT  150.0 404.7 152.7 405.9 ;
        RECT  143.7 419.4 155.1 420.6 ;
        RECT  144.9 417.3 146.1 419.4 ;
        RECT  147.9 417.3 149.1 418.5 ;
        RECT  150.9 417.3 152.1 418.5 ;
        RECT  153.9 417.3 155.1 419.4 ;
        RECT  147.6 416.4 148.8 417.3 ;
        RECT  144.9 410.7 146.1 416.4 ;
        RECT  147.6 415.2 150.0 416.4 ;
        RECT  147.6 411.9 148.8 415.2 ;
        RECT  151.2 413.7 152.4 417.3 ;
        RECT  150.6 412.5 152.4 413.7 ;
        RECT  151.2 411.9 152.4 412.5 ;
        RECT  147.3 410.7 148.5 411.9 ;
        RECT  151.5 410.7 152.7 411.9 ;
        RECT  153.9 410.7 155.1 416.4 ;
        RECT  149.4 409.2 150.6 409.5 ;
        RECT  143.7 408.0 155.1 409.2 ;
        RECT  145.8 405.9 148.5 407.1 ;
        RECT  150.0 405.9 152.7 407.1 ;
        RECT  143.7 420.6 155.1 421.8 ;
        RECT  144.9 421.8 146.1 423.9 ;
        RECT  147.9 422.7 149.1 423.9 ;
        RECT  150.9 422.7 152.1 423.9 ;
        RECT  153.9 421.8 155.1 423.9 ;
        RECT  147.6 423.9 148.8 424.8 ;
        RECT  144.9 424.8 146.1 430.5 ;
        RECT  147.6 424.8 150.0 426.0 ;
        RECT  147.6 426.0 148.8 429.3 ;
        RECT  151.2 423.9 152.4 427.5 ;
        RECT  150.6 427.5 152.4 428.7 ;
        RECT  151.2 428.7 152.4 429.3 ;
        RECT  147.3 429.3 148.5 430.5 ;
        RECT  151.5 429.3 152.7 430.5 ;
        RECT  153.9 424.8 155.1 430.5 ;
        RECT  149.4 431.7 150.6 432.0 ;
        RECT  143.7 432.0 155.1 433.2 ;
        RECT  145.8 434.1 148.5 435.3 ;
        RECT  150.0 434.1 152.7 435.3 ;
        RECT  123.9 458.4 154.5 459.3 ;
        RECT  123.9 446.4 154.5 447.3 ;
        RECT  123.9 446.4 134.1 447.3 ;
        RECT  123.9 458.4 134.1 459.3 ;
        RECT  129.3 450.9 130.2 459.3 ;
        RECT  126.9 442.5 128.1 443.7 ;
        RECT  129.3 442.5 130.5 443.7 ;
        RECT  126.9 450.9 128.1 452.1 ;
        RECT  129.3 450.9 130.5 452.1 ;
        RECT  129.3 450.9 130.5 452.1 ;
        RECT  131.7 450.9 132.9 452.1 ;
        RECT  127.8 446.4 129.0 447.6 ;
        RECT  129.3 456.3 130.5 457.5 ;
        RECT  126.9 450.9 128.1 452.1 ;
        RECT  131.7 450.9 132.9 452.1 ;
        RECT  126.9 442.5 128.1 443.7 ;
        RECT  129.3 442.5 130.5 443.7 ;
        RECT  134.1 446.4 144.3 447.3 ;
        RECT  134.1 458.4 144.3 459.3 ;
        RECT  139.5 450.9 140.4 459.3 ;
        RECT  137.1 442.5 138.3 443.7 ;
        RECT  139.5 442.5 140.7 443.7 ;
        RECT  137.1 450.9 138.3 452.1 ;
        RECT  139.5 450.9 140.7 452.1 ;
        RECT  139.5 450.9 140.7 452.1 ;
        RECT  141.9 450.9 143.1 452.1 ;
        RECT  138.0 446.4 139.2 447.6 ;
        RECT  139.5 456.3 140.7 457.5 ;
        RECT  137.1 450.9 138.3 452.1 ;
        RECT  141.9 450.9 143.1 452.1 ;
        RECT  137.1 442.5 138.3 443.7 ;
        RECT  139.5 442.5 140.7 443.7 ;
        RECT  144.3 446.4 154.5 447.3 ;
        RECT  144.3 458.4 154.5 459.3 ;
        RECT  149.7 450.9 150.6 459.3 ;
        RECT  147.3 442.5 148.5 443.7 ;
        RECT  149.7 442.5 150.9 443.7 ;
        RECT  147.3 450.9 148.5 452.1 ;
        RECT  149.7 450.9 150.9 452.1 ;
        RECT  149.7 450.9 150.9 452.1 ;
        RECT  152.1 450.9 153.3 452.1 ;
        RECT  148.2 446.4 149.4 447.6 ;
        RECT  149.7 456.3 150.9 457.5 ;
        RECT  147.3 450.9 148.5 452.1 ;
        RECT  152.1 450.9 153.3 452.1 ;
        RECT  147.3 442.5 148.5 443.7 ;
        RECT  149.7 442.5 150.9 443.7 ;
        RECT  123.9 168.75 154.5 169.65 ;
        RECT  123.9 193.95 154.5 194.85 ;
        RECT  123.9 196.05 154.5 196.95 ;
        RECT  123.3 195.9 134.7 197.1 ;
        RECT  123.3 193.8 134.7 195.0 ;
        RECT  128.7 190.2 129.9 192.9 ;
        RECT  131.1 190.2 132.3 193.8 ;
        RECT  133.5 192.6 134.7 193.8 ;
        RECT  128.7 186.3 129.6 190.2 ;
        RECT  126.0 171.9 127.2 186.3 ;
        RECT  128.4 183.6 129.6 186.3 ;
        RECT  130.8 182.7 132.0 186.3 ;
        RECT  130.8 181.5 132.9 182.7 ;
        RECT  128.4 174.6 129.6 180.0 ;
        RECT  130.8 174.6 132.0 181.5 ;
        RECT  128.4 173.7 129.3 174.6 ;
        RECT  128.4 172.8 130.2 173.7 ;
        RECT  126.0 170.7 127.8 171.9 ;
        RECT  129.3 171.0 130.2 172.8 ;
        RECT  129.3 169.8 130.5 171.0 ;
        RECT  123.3 168.6 134.7 169.8 ;
        RECT  126.6 167.4 127.8 167.7 ;
        RECT  125.7 166.5 127.8 167.4 ;
        RECT  132.6 166.5 134.1 167.7 ;
        RECT  125.7 164.4 126.6 166.5 ;
        RECT  127.8 164.4 129.0 165.6 ;
        RECT  125.7 158.1 126.9 164.4 ;
        RECT  124.8 157.2 126.9 158.1 ;
        RECT  128.1 157.2 129.3 164.4 ;
        RECT  130.5 157.2 131.7 165.6 ;
        RECT  133.2 164.4 134.1 166.5 ;
        RECT  132.9 157.2 134.1 164.4 ;
        RECT  124.8 154.5 126.0 157.2 ;
        RECT  133.5 195.9 144.9 197.1 ;
        RECT  133.5 193.8 144.9 195.0 ;
        RECT  138.9 190.2 140.1 192.9 ;
        RECT  141.3 190.2 142.5 193.8 ;
        RECT  143.7 192.6 144.9 193.8 ;
        RECT  138.9 186.3 139.8 190.2 ;
        RECT  136.2 171.9 137.4 186.3 ;
        RECT  138.6 183.6 139.8 186.3 ;
        RECT  141.0 182.7 142.2 186.3 ;
        RECT  141.0 181.5 143.1 182.7 ;
        RECT  138.6 174.6 139.8 180.0 ;
        RECT  141.0 174.6 142.2 181.5 ;
        RECT  138.6 173.7 139.5 174.6 ;
        RECT  138.6 172.8 140.4 173.7 ;
        RECT  136.2 170.7 138.0 171.9 ;
        RECT  139.5 171.0 140.4 172.8 ;
        RECT  139.5 169.8 140.7 171.0 ;
        RECT  133.5 168.6 144.9 169.8 ;
        RECT  136.8 167.4 138.0 167.7 ;
        RECT  135.9 166.5 138.0 167.4 ;
        RECT  142.8 166.5 144.3 167.7 ;
        RECT  135.9 164.4 136.8 166.5 ;
        RECT  138.0 164.4 139.2 165.6 ;
        RECT  135.9 158.1 137.1 164.4 ;
        RECT  135.0 157.2 137.1 158.1 ;
        RECT  138.3 157.2 139.5 164.4 ;
        RECT  140.7 157.2 141.9 165.6 ;
        RECT  143.4 164.4 144.3 166.5 ;
        RECT  143.1 157.2 144.3 164.4 ;
        RECT  135.0 154.5 136.2 157.2 ;
        RECT  143.7 195.9 155.1 197.1 ;
        RECT  143.7 193.8 155.1 195.0 ;
        RECT  149.1 190.2 150.3 192.9 ;
        RECT  151.5 190.2 152.7 193.8 ;
        RECT  153.9 192.6 155.1 193.8 ;
        RECT  149.1 186.3 150.0 190.2 ;
        RECT  146.4 171.9 147.6 186.3 ;
        RECT  148.8 183.6 150.0 186.3 ;
        RECT  151.2 182.7 152.4 186.3 ;
        RECT  151.2 181.5 153.3 182.7 ;
        RECT  148.8 174.6 150.0 180.0 ;
        RECT  151.2 174.6 152.4 181.5 ;
        RECT  148.8 173.7 149.7 174.6 ;
        RECT  148.8 172.8 150.6 173.7 ;
        RECT  146.4 170.7 148.2 171.9 ;
        RECT  149.7 171.0 150.6 172.8 ;
        RECT  149.7 169.8 150.9 171.0 ;
        RECT  143.7 168.6 155.1 169.8 ;
        RECT  147.0 167.4 148.2 167.7 ;
        RECT  146.1 166.5 148.2 167.4 ;
        RECT  153.0 166.5 154.5 167.7 ;
        RECT  146.1 164.4 147.0 166.5 ;
        RECT  148.2 164.4 149.4 165.6 ;
        RECT  146.1 158.1 147.3 164.4 ;
        RECT  145.2 157.2 147.3 158.1 ;
        RECT  148.5 157.2 149.7 164.4 ;
        RECT  150.9 157.2 152.1 165.6 ;
        RECT  153.6 164.4 154.5 166.5 ;
        RECT  153.3 157.2 154.5 164.4 ;
        RECT  145.2 154.5 146.4 157.2 ;
        RECT  123.9 97.95 154.5 98.85 ;
        RECT  123.9 100.05 154.5 100.95 ;
        RECT  123.9 95.85 154.5 96.75 ;
        RECT  125.4 147.9 126.6 149.1 ;
        RECT  125.4 147.3 126.3 147.9 ;
        RECT  125.1 143.7 126.3 147.3 ;
        RECT  127.5 143.7 128.7 147.3 ;
        RECT  129.9 143.7 131.1 148.5 ;
        RECT  132.3 144.9 133.8 146.1 ;
        RECT  127.8 141.3 128.7 143.7 ;
        RECT  125.1 128.1 126.3 140.7 ;
        RECT  127.8 140.1 132.0 141.3 ;
        RECT  127.2 137.7 132.0 138.9 ;
        RECT  127.5 133.8 128.7 137.7 ;
        RECT  129.9 133.2 131.1 135.0 ;
        RECT  132.9 133.2 133.8 144.9 ;
        RECT  129.9 132.0 133.8 133.2 ;
        RECT  127.5 127.2 128.7 130.2 ;
        RECT  129.9 128.1 131.1 132.0 ;
        RECT  123.9 126.0 134.7 127.2 ;
        RECT  125.4 121.8 126.6 124.8 ;
        RECT  127.8 122.7 129.0 126.0 ;
        RECT  130.2 121.8 131.4 124.8 ;
        RECT  125.4 120.9 131.4 121.8 ;
        RECT  125.4 115.2 126.6 120.9 ;
        RECT  130.2 120.6 131.4 120.9 ;
        RECT  130.2 119.4 132.0 120.6 ;
        RECT  127.8 115.2 129.0 117.3 ;
        RECT  130.2 116.4 131.4 117.3 ;
        RECT  130.2 115.2 134.1 116.4 ;
        RECT  130.8 113.1 133.2 114.3 ;
        RECT  124.8 111.9 126.0 113.1 ;
        RECT  125.1 109.8 126.0 111.9 ;
        RECT  124.8 105.9 126.0 109.8 ;
        RECT  127.2 107.7 128.4 109.8 ;
        RECT  129.6 107.7 130.8 111.0 ;
        RECT  124.8 105.0 128.4 105.9 ;
        RECT  124.8 101.1 126.0 104.1 ;
        RECT  127.2 102.0 128.4 105.0 ;
        RECT  129.6 101.1 130.8 104.1 ;
        RECT  132.0 102.0 133.2 113.1 ;
        RECT  123.9 99.9 134.7 101.1 ;
        RECT  123.9 97.8 134.7 99.0 ;
        RECT  123.9 95.7 134.7 96.9 ;
        RECT  127.5 93.6 129.9 94.8 ;
        RECT  135.6 147.9 136.8 149.1 ;
        RECT  135.6 147.3 136.5 147.9 ;
        RECT  135.3 143.7 136.5 147.3 ;
        RECT  137.7 143.7 138.9 147.3 ;
        RECT  140.1 143.7 141.3 148.5 ;
        RECT  142.5 144.9 144.0 146.1 ;
        RECT  138.0 141.3 138.9 143.7 ;
        RECT  135.3 128.1 136.5 140.7 ;
        RECT  138.0 140.1 142.2 141.3 ;
        RECT  137.4 137.7 142.2 138.9 ;
        RECT  137.7 133.8 138.9 137.7 ;
        RECT  140.1 133.2 141.3 135.0 ;
        RECT  143.1 133.2 144.0 144.9 ;
        RECT  140.1 132.0 144.0 133.2 ;
        RECT  137.7 127.2 138.9 130.2 ;
        RECT  140.1 128.1 141.3 132.0 ;
        RECT  134.1 126.0 144.9 127.2 ;
        RECT  135.6 121.8 136.8 124.8 ;
        RECT  138.0 122.7 139.2 126.0 ;
        RECT  140.4 121.8 141.6 124.8 ;
        RECT  135.6 120.9 141.6 121.8 ;
        RECT  135.6 115.2 136.8 120.9 ;
        RECT  140.4 120.6 141.6 120.9 ;
        RECT  140.4 119.4 142.2 120.6 ;
        RECT  138.0 115.2 139.2 117.3 ;
        RECT  140.4 116.4 141.6 117.3 ;
        RECT  140.4 115.2 144.3 116.4 ;
        RECT  141.0 113.1 143.4 114.3 ;
        RECT  135.0 111.9 136.2 113.1 ;
        RECT  135.3 109.8 136.2 111.9 ;
        RECT  135.0 105.9 136.2 109.8 ;
        RECT  137.4 107.7 138.6 109.8 ;
        RECT  139.8 107.7 141.0 111.0 ;
        RECT  135.0 105.0 138.6 105.9 ;
        RECT  135.0 101.1 136.2 104.1 ;
        RECT  137.4 102.0 138.6 105.0 ;
        RECT  139.8 101.1 141.0 104.1 ;
        RECT  142.2 102.0 143.4 113.1 ;
        RECT  134.1 99.9 144.9 101.1 ;
        RECT  134.1 97.8 144.9 99.0 ;
        RECT  134.1 95.7 144.9 96.9 ;
        RECT  137.7 93.6 140.1 94.8 ;
        RECT  145.8 147.9 147.0 149.1 ;
        RECT  145.8 147.3 146.7 147.9 ;
        RECT  145.5 143.7 146.7 147.3 ;
        RECT  147.9 143.7 149.1 147.3 ;
        RECT  150.3 143.7 151.5 148.5 ;
        RECT  152.7 144.9 154.2 146.1 ;
        RECT  148.2 141.3 149.1 143.7 ;
        RECT  145.5 128.1 146.7 140.7 ;
        RECT  148.2 140.1 152.4 141.3 ;
        RECT  147.6 137.7 152.4 138.9 ;
        RECT  147.9 133.8 149.1 137.7 ;
        RECT  150.3 133.2 151.5 135.0 ;
        RECT  153.3 133.2 154.2 144.9 ;
        RECT  150.3 132.0 154.2 133.2 ;
        RECT  147.9 127.2 149.1 130.2 ;
        RECT  150.3 128.1 151.5 132.0 ;
        RECT  144.3 126.0 155.1 127.2 ;
        RECT  145.8 121.8 147.0 124.8 ;
        RECT  148.2 122.7 149.4 126.0 ;
        RECT  150.6 121.8 151.8 124.8 ;
        RECT  145.8 120.9 151.8 121.8 ;
        RECT  145.8 115.2 147.0 120.9 ;
        RECT  150.6 120.6 151.8 120.9 ;
        RECT  150.6 119.4 152.4 120.6 ;
        RECT  148.2 115.2 149.4 117.3 ;
        RECT  150.6 116.4 151.8 117.3 ;
        RECT  150.6 115.2 154.5 116.4 ;
        RECT  151.2 113.1 153.6 114.3 ;
        RECT  145.2 111.9 146.4 113.1 ;
        RECT  145.5 109.8 146.4 111.9 ;
        RECT  145.2 105.9 146.4 109.8 ;
        RECT  147.6 107.7 148.8 109.8 ;
        RECT  150.0 107.7 151.2 111.0 ;
        RECT  145.2 105.0 148.8 105.9 ;
        RECT  145.2 101.1 146.4 104.1 ;
        RECT  147.6 102.0 148.8 105.0 ;
        RECT  150.0 101.1 151.2 104.1 ;
        RECT  152.4 102.0 153.6 113.1 ;
        RECT  144.3 99.9 155.1 101.1 ;
        RECT  144.3 97.8 155.1 99.0 ;
        RECT  144.3 95.7 155.1 96.9 ;
        RECT  147.9 93.6 150.3 94.8 ;
        RECT  123.9 32.85 154.5 33.75 ;
        RECT  123.9 87.3 154.5 88.2 ;
        RECT  123.3 87.3 134.7 88.2 ;
        RECT  123.3 84.0 124.5 87.3 ;
        RECT  125.7 85.5 132.3 86.4 ;
        RECT  125.7 85.2 128.7 85.5 ;
        RECT  131.1 85.2 132.3 85.5 ;
        RECT  123.3 82.8 127.5 84.0 ;
        RECT  131.1 82.8 134.7 84.0 ;
        RECT  123.3 79.2 124.5 82.8 ;
        RECT  128.7 81.9 129.9 82.8 ;
        RECT  128.7 81.6 131.1 81.9 ;
        RECT  125.7 80.7 132.3 81.6 ;
        RECT  125.7 80.4 127.5 80.7 ;
        RECT  131.1 80.4 132.3 80.7 ;
        RECT  123.3 78.0 127.5 79.2 ;
        RECT  123.3 64.2 124.5 78.0 ;
        RECT  129.0 77.4 130.2 79.8 ;
        RECT  133.8 79.2 134.7 82.8 ;
        RECT  131.1 78.0 134.7 79.2 ;
        RECT  133.5 76.8 134.7 78.0 ;
        RECT  125.7 74.4 126.9 75.6 ;
        RECT  127.8 75.3 130.2 76.5 ;
        RECT  125.7 73.5 132.3 74.4 ;
        RECT  125.7 73.2 127.5 73.5 ;
        RECT  131.1 73.2 132.3 73.5 ;
        RECT  125.7 71.1 132.3 72.0 ;
        RECT  125.7 70.8 127.5 71.1 ;
        RECT  129.9 70.8 132.3 71.1 ;
        RECT  125.7 68.7 132.3 69.6 ;
        RECT  125.7 68.4 127.5 68.7 ;
        RECT  129.9 68.4 132.3 68.7 ;
        RECT  128.7 66.6 129.9 67.5 ;
        RECT  125.7 65.7 132.3 66.6 ;
        RECT  125.7 65.4 128.7 65.7 ;
        RECT  131.1 65.4 132.3 65.7 ;
        RECT  123.3 63.0 127.5 64.2 ;
        RECT  123.3 58.5 124.5 63.0 ;
        RECT  128.4 62.1 129.6 64.5 ;
        RECT  133.8 64.2 134.7 76.8 ;
        RECT  131.1 63.0 134.7 64.2 ;
        RECT  125.7 60.9 126.9 62.1 ;
        RECT  125.7 60.0 132.3 60.9 ;
        RECT  125.7 59.7 127.5 60.0 ;
        RECT  131.1 59.7 132.3 60.0 ;
        RECT  133.8 58.5 134.7 63.0 ;
        RECT  123.3 57.3 127.5 58.5 ;
        RECT  123.3 53.7 124.5 57.3 ;
        RECT  129.0 56.4 130.2 57.6 ;
        RECT  131.1 57.3 134.7 58.5 ;
        RECT  125.7 56.1 131.1 56.4 ;
        RECT  125.7 55.5 132.3 56.1 ;
        RECT  125.7 54.9 127.5 55.5 ;
        RECT  129.9 55.2 132.3 55.5 ;
        RECT  131.1 54.9 132.3 55.2 ;
        RECT  123.3 52.5 127.5 53.7 ;
        RECT  123.3 37.5 124.5 52.5 ;
        RECT  129.0 51.9 130.2 54.3 ;
        RECT  133.8 53.7 134.7 57.3 ;
        RECT  131.1 52.5 134.7 53.7 ;
        RECT  133.5 51.3 134.7 52.5 ;
        RECT  125.7 48.0 126.9 49.2 ;
        RECT  127.8 48.9 130.2 50.1 ;
        RECT  125.7 47.1 132.3 48.0 ;
        RECT  125.7 46.8 127.5 47.1 ;
        RECT  131.1 46.8 132.3 47.1 ;
        RECT  125.7 44.7 132.3 45.6 ;
        RECT  125.7 44.4 127.5 44.7 ;
        RECT  129.9 44.4 132.3 44.7 ;
        RECT  125.7 42.3 132.3 43.2 ;
        RECT  125.7 42.0 127.5 42.3 ;
        RECT  129.9 42.0 132.3 42.3 ;
        RECT  128.7 40.2 129.9 41.1 ;
        RECT  125.7 39.3 132.3 40.2 ;
        RECT  125.7 39.0 128.7 39.3 ;
        RECT  131.1 39.0 132.3 39.3 ;
        RECT  133.8 37.8 134.7 51.3 ;
        RECT  125.7 37.5 127.5 37.8 ;
        RECT  123.3 36.6 127.5 37.5 ;
        RECT  131.1 36.9 134.7 37.8 ;
        RECT  131.1 36.6 132.3 36.9 ;
        RECT  126.3 35.1 127.5 36.6 ;
        RECT  128.4 34.2 129.6 35.1 ;
        RECT  123.3 33.3 134.7 34.2 ;
        RECT  133.5 87.3 144.9 88.2 ;
        RECT  143.7 84.0 144.9 87.3 ;
        RECT  135.9 85.5 142.5 86.4 ;
        RECT  139.5 85.2 142.5 85.5 ;
        RECT  135.9 85.2 137.1 85.5 ;
        RECT  140.7 82.8 144.9 84.0 ;
        RECT  133.5 82.8 137.1 84.0 ;
        RECT  143.7 79.2 144.9 82.8 ;
        RECT  138.3 81.9 139.5 82.8 ;
        RECT  137.1 81.6 139.5 81.9 ;
        RECT  135.9 80.7 142.5 81.6 ;
        RECT  140.7 80.4 142.5 80.7 ;
        RECT  135.9 80.4 137.1 80.7 ;
        RECT  140.7 78.0 144.9 79.2 ;
        RECT  143.7 64.2 144.9 78.0 ;
        RECT  138.0 77.4 139.2 79.8 ;
        RECT  133.5 79.2 134.4 82.8 ;
        RECT  133.5 78.0 137.1 79.2 ;
        RECT  133.5 76.8 134.7 78.0 ;
        RECT  141.3 74.4 142.5 75.6 ;
        RECT  138.0 75.3 140.4 76.5 ;
        RECT  135.9 73.5 142.5 74.4 ;
        RECT  140.7 73.2 142.5 73.5 ;
        RECT  135.9 73.2 137.1 73.5 ;
        RECT  135.9 71.1 142.5 72.0 ;
        RECT  140.7 70.8 142.5 71.1 ;
        RECT  135.9 70.8 138.3 71.1 ;
        RECT  135.9 68.7 142.5 69.6 ;
        RECT  140.7 68.4 142.5 68.7 ;
        RECT  135.9 68.4 138.3 68.7 ;
        RECT  138.3 66.6 139.5 67.5 ;
        RECT  135.9 65.7 142.5 66.6 ;
        RECT  139.5 65.4 142.5 65.7 ;
        RECT  135.9 65.4 137.1 65.7 ;
        RECT  140.7 63.0 144.9 64.2 ;
        RECT  143.7 58.5 144.9 63.0 ;
        RECT  138.6 62.1 139.8 64.5 ;
        RECT  133.5 64.2 134.4 76.8 ;
        RECT  133.5 63.0 137.1 64.2 ;
        RECT  141.3 60.9 142.5 62.1 ;
        RECT  135.9 60.0 142.5 60.9 ;
        RECT  140.7 59.7 142.5 60.0 ;
        RECT  135.9 59.7 137.1 60.0 ;
        RECT  133.5 58.5 134.4 63.0 ;
        RECT  140.7 57.3 144.9 58.5 ;
        RECT  143.7 53.7 144.9 57.3 ;
        RECT  138.0 56.4 139.2 57.6 ;
        RECT  133.5 57.3 137.1 58.5 ;
        RECT  137.1 56.1 142.5 56.4 ;
        RECT  135.9 55.5 142.5 56.1 ;
        RECT  140.7 54.9 142.5 55.5 ;
        RECT  135.9 55.2 138.3 55.5 ;
        RECT  135.9 54.9 137.1 55.2 ;
        RECT  140.7 52.5 144.9 53.7 ;
        RECT  143.7 37.5 144.9 52.5 ;
        RECT  138.0 51.9 139.2 54.3 ;
        RECT  133.5 53.7 134.4 57.3 ;
        RECT  133.5 52.5 137.1 53.7 ;
        RECT  133.5 51.3 134.7 52.5 ;
        RECT  141.3 48.0 142.5 49.2 ;
        RECT  138.0 48.9 140.4 50.1 ;
        RECT  135.9 47.1 142.5 48.0 ;
        RECT  140.7 46.8 142.5 47.1 ;
        RECT  135.9 46.8 137.1 47.1 ;
        RECT  135.9 44.7 142.5 45.6 ;
        RECT  140.7 44.4 142.5 44.7 ;
        RECT  135.9 44.4 138.3 44.7 ;
        RECT  135.9 42.3 142.5 43.2 ;
        RECT  140.7 42.0 142.5 42.3 ;
        RECT  135.9 42.0 138.3 42.3 ;
        RECT  138.3 40.2 139.5 41.1 ;
        RECT  135.9 39.3 142.5 40.2 ;
        RECT  139.5 39.0 142.5 39.3 ;
        RECT  135.9 39.0 137.1 39.3 ;
        RECT  133.5 37.8 134.4 51.3 ;
        RECT  140.7 37.5 142.5 37.8 ;
        RECT  140.7 36.6 144.9 37.5 ;
        RECT  133.5 36.9 137.1 37.8 ;
        RECT  135.9 36.6 137.1 36.9 ;
        RECT  140.7 35.1 141.9 36.6 ;
        RECT  138.6 34.2 139.8 35.1 ;
        RECT  133.5 33.3 144.9 34.2 ;
        RECT  143.7 87.3 155.1 88.2 ;
        RECT  143.7 84.0 144.9 87.3 ;
        RECT  146.1 85.5 152.7 86.4 ;
        RECT  146.1 85.2 149.1 85.5 ;
        RECT  151.5 85.2 152.7 85.5 ;
        RECT  143.7 82.8 147.9 84.0 ;
        RECT  151.5 82.8 155.1 84.0 ;
        RECT  143.7 79.2 144.9 82.8 ;
        RECT  149.1 81.9 150.3 82.8 ;
        RECT  149.1 81.6 151.5 81.9 ;
        RECT  146.1 80.7 152.7 81.6 ;
        RECT  146.1 80.4 147.9 80.7 ;
        RECT  151.5 80.4 152.7 80.7 ;
        RECT  143.7 78.0 147.9 79.2 ;
        RECT  143.7 64.2 144.9 78.0 ;
        RECT  149.4 77.4 150.6 79.8 ;
        RECT  154.2 79.2 155.1 82.8 ;
        RECT  151.5 78.0 155.1 79.2 ;
        RECT  153.9 76.8 155.1 78.0 ;
        RECT  146.1 74.4 147.3 75.6 ;
        RECT  148.2 75.3 150.6 76.5 ;
        RECT  146.1 73.5 152.7 74.4 ;
        RECT  146.1 73.2 147.9 73.5 ;
        RECT  151.5 73.2 152.7 73.5 ;
        RECT  146.1 71.1 152.7 72.0 ;
        RECT  146.1 70.8 147.9 71.1 ;
        RECT  150.3 70.8 152.7 71.1 ;
        RECT  146.1 68.7 152.7 69.6 ;
        RECT  146.1 68.4 147.9 68.7 ;
        RECT  150.3 68.4 152.7 68.7 ;
        RECT  149.1 66.6 150.3 67.5 ;
        RECT  146.1 65.7 152.7 66.6 ;
        RECT  146.1 65.4 149.1 65.7 ;
        RECT  151.5 65.4 152.7 65.7 ;
        RECT  143.7 63.0 147.9 64.2 ;
        RECT  143.7 58.5 144.9 63.0 ;
        RECT  148.8 62.1 150.0 64.5 ;
        RECT  154.2 64.2 155.1 76.8 ;
        RECT  151.5 63.0 155.1 64.2 ;
        RECT  146.1 60.9 147.3 62.1 ;
        RECT  146.1 60.0 152.7 60.9 ;
        RECT  146.1 59.7 147.9 60.0 ;
        RECT  151.5 59.7 152.7 60.0 ;
        RECT  154.2 58.5 155.1 63.0 ;
        RECT  143.7 57.3 147.9 58.5 ;
        RECT  143.7 53.7 144.9 57.3 ;
        RECT  149.4 56.4 150.6 57.6 ;
        RECT  151.5 57.3 155.1 58.5 ;
        RECT  146.1 56.1 151.5 56.4 ;
        RECT  146.1 55.5 152.7 56.1 ;
        RECT  146.1 54.9 147.9 55.5 ;
        RECT  150.3 55.2 152.7 55.5 ;
        RECT  151.5 54.9 152.7 55.2 ;
        RECT  143.7 52.5 147.9 53.7 ;
        RECT  143.7 37.5 144.9 52.5 ;
        RECT  149.4 51.9 150.6 54.3 ;
        RECT  154.2 53.7 155.1 57.3 ;
        RECT  151.5 52.5 155.1 53.7 ;
        RECT  153.9 51.3 155.1 52.5 ;
        RECT  146.1 48.0 147.3 49.2 ;
        RECT  148.2 48.9 150.6 50.1 ;
        RECT  146.1 47.1 152.7 48.0 ;
        RECT  146.1 46.8 147.9 47.1 ;
        RECT  151.5 46.8 152.7 47.1 ;
        RECT  146.1 44.7 152.7 45.6 ;
        RECT  146.1 44.4 147.9 44.7 ;
        RECT  150.3 44.4 152.7 44.7 ;
        RECT  146.1 42.3 152.7 43.2 ;
        RECT  146.1 42.0 147.9 42.3 ;
        RECT  150.3 42.0 152.7 42.3 ;
        RECT  149.1 40.2 150.3 41.1 ;
        RECT  146.1 39.3 152.7 40.2 ;
        RECT  146.1 39.0 149.1 39.3 ;
        RECT  151.5 39.0 152.7 39.3 ;
        RECT  154.2 37.8 155.1 51.3 ;
        RECT  146.1 37.5 147.9 37.8 ;
        RECT  143.7 36.6 147.9 37.5 ;
        RECT  151.5 36.9 155.1 37.8 ;
        RECT  151.5 36.6 152.7 36.9 ;
        RECT  146.7 35.1 147.9 36.6 ;
        RECT  148.8 34.2 150.0 35.1 ;
        RECT  143.7 33.3 155.1 34.2 ;
        RECT  123.9 26.25 154.5 27.15 ;
        RECT  123.9 28.65 154.5 29.55 ;
        RECT  123.9 10.35 154.5 11.25 ;
        RECT  123.9 50.4 134.7 51.6 ;
        RECT  124.8 46.8 126.3 49.2 ;
        RECT  127.5 46.8 128.7 50.4 ;
        RECT  129.9 46.8 131.1 49.2 ;
        RECT  132.3 46.8 133.5 49.2 ;
        RECT  124.8 43.5 125.7 46.8 ;
        RECT  126.6 44.7 127.8 45.9 ;
        RECT  124.8 42.3 129.9 43.5 ;
        RECT  132.6 42.3 133.5 46.8 ;
        RECT  124.8 40.2 125.7 42.3 ;
        RECT  131.4 41.1 133.5 42.3 ;
        RECT  132.6 40.2 133.5 41.1 ;
        RECT  124.8 39.0 126.3 40.2 ;
        RECT  127.5 37.8 128.7 40.2 ;
        RECT  129.9 39.0 131.1 40.2 ;
        RECT  132.3 39.0 133.5 40.2 ;
        RECT  123.9 36.6 134.7 37.8 ;
        RECT  123.9 34.5 134.7 35.7 ;
        RECT  123.9 32.1 134.7 33.3 ;
        RECT  133.5 50.4 144.3 51.6 ;
        RECT  141.9 46.8 143.4 49.2 ;
        RECT  139.5 46.8 140.7 50.4 ;
        RECT  137.1 46.8 138.3 49.2 ;
        RECT  134.7 46.8 135.9 49.2 ;
        RECT  142.5 43.5 143.4 46.8 ;
        RECT  140.4 44.7 141.6 45.9 ;
        RECT  138.3 42.3 143.4 43.5 ;
        RECT  134.7 42.3 135.6 46.8 ;
        RECT  142.5 40.2 143.4 42.3 ;
        RECT  134.7 41.1 136.8 42.3 ;
        RECT  134.7 40.2 135.6 41.1 ;
        RECT  141.9 39.0 143.4 40.2 ;
        RECT  139.5 37.8 140.7 40.2 ;
        RECT  137.1 39.0 138.3 40.2 ;
        RECT  134.7 39.0 135.9 40.2 ;
        RECT  133.5 36.6 144.3 37.8 ;
        RECT  133.5 34.5 144.3 35.7 ;
        RECT  133.5 32.1 144.3 33.3 ;
        RECT  144.3 50.4 155.1 51.6 ;
        RECT  145.2 46.8 146.7 49.2 ;
        RECT  147.9 46.8 149.1 50.4 ;
        RECT  150.3 46.8 151.5 49.2 ;
        RECT  152.7 46.8 153.9 49.2 ;
        RECT  145.2 43.5 146.1 46.8 ;
        RECT  147.0 44.7 148.2 45.9 ;
        RECT  145.2 42.3 150.3 43.5 ;
        RECT  153.0 42.3 153.9 46.8 ;
        RECT  145.2 40.2 146.1 42.3 ;
        RECT  151.8 41.1 153.9 42.3 ;
        RECT  153.0 40.2 153.9 41.1 ;
        RECT  145.2 39.0 146.7 40.2 ;
        RECT  147.9 37.8 149.1 40.2 ;
        RECT  150.3 39.0 151.5 40.2 ;
        RECT  152.7 39.0 153.9 40.2 ;
        RECT  144.3 36.6 155.1 37.8 ;
        RECT  144.3 34.5 155.1 35.7 ;
        RECT  144.3 32.1 155.1 33.3 ;
        RECT  41.4 206.4 42.3 207.3 ;
        RECT  41.4 222.3 42.3 223.2 ;
        RECT  41.4 235.8 42.3 236.7 ;
        RECT  41.4 251.7 42.3 252.6 ;
        RECT  41.4 265.2 42.3 266.1 ;
        RECT  41.4 281.1 42.3 282.0 ;
        RECT  41.4 294.6 42.3 295.5 ;
        RECT  41.4 310.5 42.3 311.4 ;
        RECT  41.4 324.0 42.3 324.9 ;
        RECT  41.4 339.9 42.3 340.8 ;
        RECT  41.4 353.4 42.3 354.3 ;
        RECT  41.4 369.3 42.3 370.2 ;
        RECT  41.4 382.8 42.3 383.7 ;
        RECT  41.4 398.7 42.3 399.6 ;
        RECT  41.4 412.2 42.3 413.1 ;
        RECT  41.4 428.1 42.3 429.0 ;
        RECT  12.6 88.8 29.4 89.7 ;
        RECT  14.7 104.7 29.4 105.6 ;
        RECT  16.8 118.2 29.4 119.1 ;
        RECT  18.9 134.1 29.4 135.0 ;
        RECT  21.0 147.6 29.4 148.5 ;
        RECT  23.1 163.5 29.4 164.4 ;
        RECT  25.2 177.0 29.4 177.9 ;
        RECT  27.3 192.9 29.4 193.8 ;
        RECT  12.6 208.8 29.4 209.7 ;
        RECT  21.0 205.5 29.4 206.4 ;
        RECT  12.6 219.9 29.4 220.8 ;
        RECT  23.1 223.2 29.4 224.1 ;
        RECT  12.6 238.2 29.4 239.1 ;
        RECT  25.2 234.9 29.4 235.8 ;
        RECT  12.6 249.3 29.4 250.2 ;
        RECT  27.3 252.6 29.4 253.5 ;
        RECT  14.7 267.6 29.4 268.5 ;
        RECT  21.0 264.3 29.4 265.2 ;
        RECT  14.7 278.7 29.4 279.6 ;
        RECT  23.1 282.0 29.4 282.9 ;
        RECT  14.7 297.0 29.4 297.9 ;
        RECT  25.2 293.7 29.4 294.6 ;
        RECT  14.7 308.1 29.4 309.0 ;
        RECT  27.3 311.4 29.4 312.3 ;
        RECT  16.8 326.4 29.4 327.3 ;
        RECT  21.0 323.1 29.4 324.0 ;
        RECT  16.8 337.5 29.4 338.4 ;
        RECT  23.1 340.8 29.4 341.7 ;
        RECT  16.8 355.8 29.4 356.7 ;
        RECT  25.2 352.5 29.4 353.4 ;
        RECT  16.8 366.9 29.4 367.8 ;
        RECT  27.3 370.2 29.4 371.1 ;
        RECT  18.9 385.2 29.4 386.1 ;
        RECT  21.0 381.9 29.4 382.8 ;
        RECT  18.9 396.3 29.4 397.2 ;
        RECT  23.1 399.6 29.4 400.5 ;
        RECT  18.9 414.6 29.4 415.5 ;
        RECT  25.2 411.3 29.4 412.2 ;
        RECT  18.9 425.7 29.4 426.6 ;
        RECT  27.3 429.0 29.4 429.9 ;
        RECT  38.1 88.8 39.0 89.7 ;
        RECT  38.1 104.7 39.0 105.6 ;
        RECT  38.1 118.2 39.0 119.1 ;
        RECT  38.1 134.1 39.0 135.0 ;
        RECT  63.9 88.8 64.8 94.95 ;
        RECT  58.5 94.05 64.8 94.95 ;
        RECT  73.5 88.8 78.6 89.7 ;
        RECT  62.7 96.75 74.4 97.65 ;
        RECT  60.6 82.05 74.4 82.95 ;
        RECT  63.9 99.45 64.8 105.6 ;
        RECT  56.4 99.45 64.8 100.35 ;
        RECT  73.5 104.7 76.5 105.6 ;
        RECT  62.7 96.75 74.4 97.65 ;
        RECT  60.6 111.45 74.4 112.35 ;
        RECT  51.0 91.2 59.4 92.1 ;
        RECT  51.0 87.9 57.3 88.8 ;
        RECT  51.0 102.3 55.2 103.2 ;
        RECT  51.0 105.6 57.3 106.5 ;
        RECT  51.0 120.6 59.4 121.5 ;
        RECT  51.0 117.3 53.1 118.2 ;
        RECT  51.0 131.7 55.2 132.6 ;
        RECT  51.0 131.7 78.6 132.6 ;
        RECT  51.0 135.0 53.1 135.9 ;
        RECT  51.0 135.0 76.5 135.9 ;
        RECT  51.0 82.05 61.5 82.95 ;
        RECT  51.0 96.75 63.6 97.65 ;
        RECT  51.0 111.45 61.5 112.35 ;
        RECT  51.0 126.15 63.6 127.05 ;
        RECT  51.0 140.85 61.5 141.75 ;
        RECT  60.6 138.6 61.5 140.85 ;
        RECT  64.8 82.05 74.4 82.95 ;
        RECT  64.8 67.35 74.4 68.25 ;
        RECT  66.6 68.25 67.8 70.65 ;
        RECT  66.6 80.25 67.8 82.05 ;
        RECT  71.4 81.15 72.6 82.05 ;
        RECT  71.4 68.25 72.6 69.45 ;
        RECT  69.0 70.5 70.2 79.95 ;
        RECT  72.3 75.3 74.4 76.2 ;
        RECT  64.8 75.3 69.0 76.2 ;
        RECT  71.4 78.75 72.6 79.95 ;
        RECT  69.0 78.75 70.2 79.95 ;
        RECT  71.4 69.45 72.6 70.65 ;
        RECT  69.0 69.45 70.2 70.65 ;
        RECT  66.6 69.45 67.8 70.65 ;
        RECT  66.6 79.95 67.8 81.15 ;
        RECT  71.1 75.15 72.3 76.35 ;
        RECT  64.8 111.45 74.4 112.35 ;
        RECT  64.8 126.15 74.4 127.05 ;
        RECT  66.6 123.75 67.8 126.15 ;
        RECT  66.6 112.35 67.8 114.15 ;
        RECT  71.4 112.35 72.6 113.25 ;
        RECT  71.4 124.95 72.6 126.15 ;
        RECT  69.0 114.45 70.2 123.9 ;
        RECT  72.3 118.2 74.4 119.1 ;
        RECT  64.8 118.2 69.0 119.1 ;
        RECT  71.4 116.85 72.6 118.05 ;
        RECT  69.0 116.85 70.2 118.05 ;
        RECT  71.4 117.75 72.6 118.95 ;
        RECT  69.0 117.75 70.2 118.95 ;
        RECT  66.6 122.55 67.8 123.75 ;
        RECT  66.6 112.05 67.8 113.25 ;
        RECT  71.1 116.85 72.3 118.05 ;
        RECT  29.4 82.05 39.0 82.95 ;
        RECT  29.4 67.35 39.0 68.25 ;
        RECT  31.2 68.25 32.4 70.65 ;
        RECT  31.2 80.25 32.4 82.05 ;
        RECT  36.0 81.15 37.2 82.05 ;
        RECT  36.0 68.25 37.2 69.45 ;
        RECT  33.6 70.5 34.8 79.95 ;
        RECT  36.9 75.3 39.0 76.2 ;
        RECT  29.4 75.3 33.6 76.2 ;
        RECT  36.0 78.75 37.2 79.95 ;
        RECT  33.6 78.75 34.8 79.95 ;
        RECT  36.0 69.45 37.2 70.65 ;
        RECT  33.6 69.45 34.8 70.65 ;
        RECT  31.2 69.45 32.4 70.65 ;
        RECT  31.2 79.95 32.4 81.15 ;
        RECT  35.7 75.15 36.9 76.35 ;
        RECT  29.4 111.45 39.0 112.35 ;
        RECT  29.4 126.15 39.0 127.05 ;
        RECT  31.2 123.75 32.4 126.15 ;
        RECT  31.2 112.35 32.4 114.15 ;
        RECT  36.0 112.35 37.2 113.25 ;
        RECT  36.0 124.95 37.2 126.15 ;
        RECT  33.6 114.45 34.8 123.9 ;
        RECT  36.9 118.2 39.0 119.1 ;
        RECT  29.4 118.2 33.6 119.1 ;
        RECT  36.0 116.85 37.2 118.05 ;
        RECT  33.6 116.85 34.8 118.05 ;
        RECT  36.0 117.75 37.2 118.95 ;
        RECT  33.6 117.75 34.8 118.95 ;
        RECT  31.2 122.55 32.4 123.75 ;
        RECT  31.2 112.05 32.4 113.25 ;
        RECT  35.7 116.85 36.9 118.05 ;
        RECT  29.4 111.45 39.0 112.35 ;
        RECT  29.4 96.75 39.0 97.65 ;
        RECT  31.2 97.65 32.4 100.05 ;
        RECT  31.2 109.65 32.4 111.45 ;
        RECT  36.0 110.55 37.2 111.45 ;
        RECT  36.0 97.65 37.2 98.85 ;
        RECT  33.6 99.9 34.8 109.35 ;
        RECT  36.9 104.7 39.0 105.6 ;
        RECT  29.4 104.7 33.6 105.6 ;
        RECT  36.0 108.15 37.2 109.35 ;
        RECT  33.6 108.15 34.8 109.35 ;
        RECT  36.0 98.85 37.2 100.05 ;
        RECT  33.6 98.85 34.8 100.05 ;
        RECT  31.2 98.85 32.4 100.05 ;
        RECT  31.2 109.35 32.4 110.55 ;
        RECT  35.7 104.55 36.9 105.75 ;
        RECT  29.4 140.85 39.0 141.75 ;
        RECT  29.4 155.55 39.0 156.45 ;
        RECT  31.2 153.15 32.4 155.55 ;
        RECT  31.2 141.75 32.4 143.55 ;
        RECT  36.0 141.75 37.2 142.65 ;
        RECT  36.0 154.35 37.2 155.55 ;
        RECT  33.6 143.85 34.8 153.3 ;
        RECT  36.9 147.6 39.0 148.5 ;
        RECT  29.4 147.6 33.6 148.5 ;
        RECT  36.0 146.25 37.2 147.45 ;
        RECT  33.6 146.25 34.8 147.45 ;
        RECT  36.0 147.15 37.2 148.35 ;
        RECT  33.6 147.15 34.8 148.35 ;
        RECT  31.2 151.95 32.4 153.15 ;
        RECT  31.2 141.45 32.4 142.65 ;
        RECT  35.7 146.25 36.9 147.45 ;
        RECT  39.0 82.05 51.0 82.95 ;
        RECT  39.0 67.35 51.0 68.25 ;
        RECT  41.1 67.8 42.0 70.65 ;
        RECT  41.1 80.1 42.0 82.5 ;
        RECT  48.15 67.8 49.05 70.65 ;
        RECT  43.35 67.8 44.25 70.65 ;
        RECT  48.15 79.65 49.05 82.5 ;
        RECT  48.9 72.9 51.0 73.8 ;
        RECT  45.9 76.2 51.0 77.1 ;
        RECT  39.0 75.3 43.35 76.2 ;
        RECT  48.0 78.45 49.2 79.65 ;
        RECT  45.6 78.45 46.8 79.65 ;
        RECT  45.6 78.45 46.8 79.65 ;
        RECT  43.2 78.45 44.4 79.65 ;
        RECT  48.0 69.45 49.2 70.65 ;
        RECT  45.6 69.45 46.8 70.65 ;
        RECT  45.6 69.45 46.8 70.65 ;
        RECT  43.2 69.45 44.4 70.65 ;
        RECT  40.8 69.45 42.0 70.65 ;
        RECT  40.8 79.65 42.0 80.85 ;
        RECT  42.9 72.9 43.8 73.8 ;
        RECT  45.9 72.9 46.8 73.8 ;
        RECT  42.9 73.35 43.8 80.85 ;
        RECT  43.35 72.9 46.35 73.8 ;
        RECT  45.9 70.65 46.8 73.35 ;
        RECT  47.7 72.9 48.9 74.1 ;
        RECT  44.7 76.2 45.9 77.4 ;
        RECT  39.0 111.45 51.0 112.35 ;
        RECT  39.0 126.15 51.0 127.05 ;
        RECT  41.1 123.75 42.0 126.6 ;
        RECT  41.1 111.9 42.0 114.3 ;
        RECT  48.15 123.75 49.05 126.6 ;
        RECT  43.35 123.75 44.25 126.6 ;
        RECT  48.15 111.9 49.05 114.75 ;
        RECT  48.9 120.6 51.0 121.5 ;
        RECT  45.9 117.3 51.0 118.2 ;
        RECT  39.0 118.2 43.35 119.1 ;
        RECT  48.0 118.35 49.2 119.55 ;
        RECT  45.6 118.35 46.8 119.55 ;
        RECT  45.6 118.35 46.8 119.55 ;
        RECT  43.2 118.35 44.4 119.55 ;
        RECT  48.0 117.75 49.2 118.95 ;
        RECT  45.6 117.75 46.8 118.95 ;
        RECT  45.6 117.75 46.8 118.95 ;
        RECT  43.2 117.75 44.4 118.95 ;
        RECT  40.8 122.55 42.0 123.75 ;
        RECT  40.8 112.35 42.0 113.55 ;
        RECT  42.9 105.6 43.8 106.5 ;
        RECT  45.9 105.6 46.8 106.5 ;
        RECT  42.9 106.05 43.8 113.55 ;
        RECT  43.35 105.6 46.35 106.5 ;
        RECT  45.9 103.35 46.8 106.05 ;
        RECT  47.7 119.1 48.9 120.3 ;
        RECT  44.7 115.8 45.9 117.0 ;
        RECT  39.0 111.45 51.0 112.35 ;
        RECT  39.0 96.75 51.0 97.65 ;
        RECT  41.1 97.2 42.0 100.05 ;
        RECT  41.1 109.5 42.0 111.9 ;
        RECT  48.15 97.2 49.05 100.05 ;
        RECT  43.35 97.2 44.25 100.05 ;
        RECT  48.15 109.05 49.05 111.9 ;
        RECT  48.9 102.3 51.0 103.2 ;
        RECT  45.9 105.6 51.0 106.5 ;
        RECT  39.0 104.7 43.35 105.6 ;
        RECT  48.0 107.85 49.2 109.05 ;
        RECT  45.6 107.85 46.8 109.05 ;
        RECT  45.6 107.85 46.8 109.05 ;
        RECT  43.2 107.85 44.4 109.05 ;
        RECT  48.0 98.85 49.2 100.05 ;
        RECT  45.6 98.85 46.8 100.05 ;
        RECT  45.6 98.85 46.8 100.05 ;
        RECT  43.2 98.85 44.4 100.05 ;
        RECT  40.8 98.85 42.0 100.05 ;
        RECT  40.8 109.05 42.0 110.25 ;
        RECT  42.9 102.3 43.8 103.2 ;
        RECT  45.9 102.3 46.8 103.2 ;
        RECT  42.9 102.75 43.8 110.25 ;
        RECT  43.35 102.3 46.35 103.2 ;
        RECT  45.9 100.05 46.8 102.75 ;
        RECT  47.7 102.3 48.9 103.5 ;
        RECT  44.7 105.6 45.9 106.8 ;
        RECT  39.0 140.85 51.0 141.75 ;
        RECT  39.0 155.55 51.0 156.45 ;
        RECT  41.1 153.15 42.0 156.0 ;
        RECT  41.1 141.3 42.0 143.7 ;
        RECT  48.15 153.15 49.05 156.0 ;
        RECT  43.35 153.15 44.25 156.0 ;
        RECT  48.15 141.3 49.05 144.15 ;
        RECT  48.9 150.0 51.0 150.9 ;
        RECT  45.9 146.7 51.0 147.6 ;
        RECT  39.0 147.6 43.35 148.5 ;
        RECT  48.0 147.75 49.2 148.95 ;
        RECT  45.6 147.75 46.8 148.95 ;
        RECT  45.6 147.75 46.8 148.95 ;
        RECT  43.2 147.75 44.4 148.95 ;
        RECT  48.0 147.15 49.2 148.35 ;
        RECT  45.6 147.15 46.8 148.35 ;
        RECT  45.6 147.15 46.8 148.35 ;
        RECT  43.2 147.15 44.4 148.35 ;
        RECT  40.8 151.95 42.0 153.15 ;
        RECT  40.8 141.75 42.0 142.95 ;
        RECT  42.9 135.0 43.8 135.9 ;
        RECT  45.9 135.0 46.8 135.9 ;
        RECT  42.9 135.45 43.8 142.95 ;
        RECT  43.35 135.0 46.35 135.9 ;
        RECT  45.9 132.75 46.8 135.45 ;
        RECT  47.7 148.5 48.9 149.7 ;
        RECT  44.7 145.2 45.9 146.4 ;
        RECT  58.2 92.85 59.4 94.05 ;
        RECT  77.4 87.6 78.6 88.8 ;
        RECT  56.1 98.25 57.3 99.45 ;
        RECT  75.3 103.5 76.5 104.7 ;
        RECT  58.2 90.0 59.4 91.2 ;
        RECT  56.1 86.7 57.3 87.9 ;
        RECT  54.0 101.1 55.2 102.3 ;
        RECT  56.1 104.4 57.3 105.6 ;
        RECT  58.2 119.4 59.4 120.6 ;
        RECT  51.9 116.1 53.1 117.3 ;
        RECT  54.0 130.5 55.2 131.7 ;
        RECT  77.4 130.5 78.6 131.7 ;
        RECT  51.9 133.8 53.1 135.0 ;
        RECT  75.3 133.8 76.5 135.0 ;
        RECT  60.3 80.85 61.5 82.05 ;
        RECT  62.4 95.55 63.6 96.75 ;
        RECT  60.3 110.25 61.5 111.45 ;
        RECT  62.4 124.95 63.6 126.15 ;
        RECT  60.3 137.4 61.5 138.6 ;
        RECT  38.1 147.6 39.0 148.5 ;
        RECT  38.1 163.5 39.0 164.4 ;
        RECT  38.1 177.0 39.0 177.9 ;
        RECT  38.1 192.9 39.0 193.8 ;
        RECT  63.9 147.6 64.8 153.75 ;
        RECT  58.5 152.85 64.8 153.75 ;
        RECT  73.5 147.6 78.6 148.5 ;
        RECT  62.7 155.55 74.4 156.45 ;
        RECT  60.6 140.85 74.4 141.75 ;
        RECT  63.9 158.25 64.8 164.4 ;
        RECT  56.4 158.25 64.8 159.15 ;
        RECT  73.5 163.5 76.5 164.4 ;
        RECT  62.7 155.55 74.4 156.45 ;
        RECT  60.6 170.25 74.4 171.15 ;
        RECT  51.0 150.0 59.4 150.9 ;
        RECT  51.0 146.7 57.3 147.6 ;
        RECT  51.0 161.1 55.2 162.0 ;
        RECT  51.0 164.4 57.3 165.3 ;
        RECT  51.0 179.4 59.4 180.3 ;
        RECT  51.0 176.1 53.1 177.0 ;
        RECT  51.0 190.5 55.2 191.4 ;
        RECT  51.0 190.5 78.6 191.4 ;
        RECT  51.0 193.8 53.1 194.7 ;
        RECT  51.0 193.8 76.5 194.7 ;
        RECT  51.0 140.85 61.5 141.75 ;
        RECT  51.0 155.55 63.6 156.45 ;
        RECT  51.0 170.25 61.5 171.15 ;
        RECT  51.0 184.95 63.6 185.85 ;
        RECT  51.0 199.65 61.5 200.55 ;
        RECT  60.6 197.4 61.5 199.65 ;
        RECT  64.8 140.85 74.4 141.75 ;
        RECT  64.8 126.15 74.4 127.05 ;
        RECT  66.6 127.05 67.8 129.45 ;
        RECT  66.6 139.05 67.8 140.85 ;
        RECT  71.4 139.95 72.6 140.85 ;
        RECT  71.4 127.05 72.6 128.25 ;
        RECT  69.0 129.3 70.2 138.75 ;
        RECT  72.3 134.1 74.4 135.0 ;
        RECT  64.8 134.1 69.0 135.0 ;
        RECT  71.4 137.55 72.6 138.75 ;
        RECT  69.0 137.55 70.2 138.75 ;
        RECT  71.4 128.25 72.6 129.45 ;
        RECT  69.0 128.25 70.2 129.45 ;
        RECT  66.6 128.25 67.8 129.45 ;
        RECT  66.6 138.75 67.8 139.95 ;
        RECT  71.1 133.95 72.3 135.15 ;
        RECT  64.8 170.25 74.4 171.15 ;
        RECT  64.8 184.95 74.4 185.85 ;
        RECT  66.6 182.55 67.8 184.95 ;
        RECT  66.6 171.15 67.8 172.95 ;
        RECT  71.4 171.15 72.6 172.05 ;
        RECT  71.4 183.75 72.6 184.95 ;
        RECT  69.0 173.25 70.2 182.7 ;
        RECT  72.3 177.0 74.4 177.9 ;
        RECT  64.8 177.0 69.0 177.9 ;
        RECT  71.4 175.65 72.6 176.85 ;
        RECT  69.0 175.65 70.2 176.85 ;
        RECT  71.4 176.55 72.6 177.75 ;
        RECT  69.0 176.55 70.2 177.75 ;
        RECT  66.6 181.35 67.8 182.55 ;
        RECT  66.6 170.85 67.8 172.05 ;
        RECT  71.1 175.65 72.3 176.85 ;
        RECT  29.4 140.85 39.0 141.75 ;
        RECT  29.4 126.15 39.0 127.05 ;
        RECT  31.2 127.05 32.4 129.45 ;
        RECT  31.2 139.05 32.4 140.85 ;
        RECT  36.0 139.95 37.2 140.85 ;
        RECT  36.0 127.05 37.2 128.25 ;
        RECT  33.6 129.3 34.8 138.75 ;
        RECT  36.9 134.1 39.0 135.0 ;
        RECT  29.4 134.1 33.6 135.0 ;
        RECT  36.0 137.55 37.2 138.75 ;
        RECT  33.6 137.55 34.8 138.75 ;
        RECT  36.0 128.25 37.2 129.45 ;
        RECT  33.6 128.25 34.8 129.45 ;
        RECT  31.2 128.25 32.4 129.45 ;
        RECT  31.2 138.75 32.4 139.95 ;
        RECT  35.7 133.95 36.9 135.15 ;
        RECT  29.4 170.25 39.0 171.15 ;
        RECT  29.4 184.95 39.0 185.85 ;
        RECT  31.2 182.55 32.4 184.95 ;
        RECT  31.2 171.15 32.4 172.95 ;
        RECT  36.0 171.15 37.2 172.05 ;
        RECT  36.0 183.75 37.2 184.95 ;
        RECT  33.6 173.25 34.8 182.7 ;
        RECT  36.9 177.0 39.0 177.9 ;
        RECT  29.4 177.0 33.6 177.9 ;
        RECT  36.0 175.65 37.2 176.85 ;
        RECT  33.6 175.65 34.8 176.85 ;
        RECT  36.0 176.55 37.2 177.75 ;
        RECT  33.6 176.55 34.8 177.75 ;
        RECT  31.2 181.35 32.4 182.55 ;
        RECT  31.2 170.85 32.4 172.05 ;
        RECT  35.7 175.65 36.9 176.85 ;
        RECT  29.4 170.25 39.0 171.15 ;
        RECT  29.4 155.55 39.0 156.45 ;
        RECT  31.2 156.45 32.4 158.85 ;
        RECT  31.2 168.45 32.4 170.25 ;
        RECT  36.0 169.35 37.2 170.25 ;
        RECT  36.0 156.45 37.2 157.65 ;
        RECT  33.6 158.7 34.8 168.15 ;
        RECT  36.9 163.5 39.0 164.4 ;
        RECT  29.4 163.5 33.6 164.4 ;
        RECT  36.0 166.95 37.2 168.15 ;
        RECT  33.6 166.95 34.8 168.15 ;
        RECT  36.0 157.65 37.2 158.85 ;
        RECT  33.6 157.65 34.8 158.85 ;
        RECT  31.2 157.65 32.4 158.85 ;
        RECT  31.2 168.15 32.4 169.35 ;
        RECT  35.7 163.35 36.9 164.55 ;
        RECT  29.4 199.65 39.0 200.55 ;
        RECT  29.4 214.35 39.0 215.25 ;
        RECT  31.2 211.95 32.4 214.35 ;
        RECT  31.2 200.55 32.4 202.35 ;
        RECT  36.0 200.55 37.2 201.45 ;
        RECT  36.0 213.15 37.2 214.35 ;
        RECT  33.6 202.65 34.8 212.1 ;
        RECT  36.9 206.4 39.0 207.3 ;
        RECT  29.4 206.4 33.6 207.3 ;
        RECT  36.0 205.05 37.2 206.25 ;
        RECT  33.6 205.05 34.8 206.25 ;
        RECT  36.0 205.95 37.2 207.15 ;
        RECT  33.6 205.95 34.8 207.15 ;
        RECT  31.2 210.75 32.4 211.95 ;
        RECT  31.2 200.25 32.4 201.45 ;
        RECT  35.7 205.05 36.9 206.25 ;
        RECT  39.0 140.85 51.0 141.75 ;
        RECT  39.0 126.15 51.0 127.05 ;
        RECT  41.1 126.6 42.0 129.45 ;
        RECT  41.1 138.9 42.0 141.3 ;
        RECT  48.15 126.6 49.05 129.45 ;
        RECT  43.35 126.6 44.25 129.45 ;
        RECT  48.15 138.45 49.05 141.3 ;
        RECT  48.9 131.7 51.0 132.6 ;
        RECT  45.9 135.0 51.0 135.9 ;
        RECT  39.0 134.1 43.35 135.0 ;
        RECT  48.0 137.25 49.2 138.45 ;
        RECT  45.6 137.25 46.8 138.45 ;
        RECT  45.6 137.25 46.8 138.45 ;
        RECT  43.2 137.25 44.4 138.45 ;
        RECT  48.0 128.25 49.2 129.45 ;
        RECT  45.6 128.25 46.8 129.45 ;
        RECT  45.6 128.25 46.8 129.45 ;
        RECT  43.2 128.25 44.4 129.45 ;
        RECT  40.8 128.25 42.0 129.45 ;
        RECT  40.8 138.45 42.0 139.65 ;
        RECT  42.9 131.7 43.8 132.6 ;
        RECT  45.9 131.7 46.8 132.6 ;
        RECT  42.9 132.15 43.8 139.65 ;
        RECT  43.35 131.7 46.35 132.6 ;
        RECT  45.9 129.45 46.8 132.15 ;
        RECT  47.7 131.7 48.9 132.9 ;
        RECT  44.7 135.0 45.9 136.2 ;
        RECT  39.0 170.25 51.0 171.15 ;
        RECT  39.0 184.95 51.0 185.85 ;
        RECT  41.1 182.55 42.0 185.4 ;
        RECT  41.1 170.7 42.0 173.1 ;
        RECT  48.15 182.55 49.05 185.4 ;
        RECT  43.35 182.55 44.25 185.4 ;
        RECT  48.15 170.7 49.05 173.55 ;
        RECT  48.9 179.4 51.0 180.3 ;
        RECT  45.9 176.1 51.0 177.0 ;
        RECT  39.0 177.0 43.35 177.9 ;
        RECT  48.0 177.15 49.2 178.35 ;
        RECT  45.6 177.15 46.8 178.35 ;
        RECT  45.6 177.15 46.8 178.35 ;
        RECT  43.2 177.15 44.4 178.35 ;
        RECT  48.0 176.55 49.2 177.75 ;
        RECT  45.6 176.55 46.8 177.75 ;
        RECT  45.6 176.55 46.8 177.75 ;
        RECT  43.2 176.55 44.4 177.75 ;
        RECT  40.8 181.35 42.0 182.55 ;
        RECT  40.8 171.15 42.0 172.35 ;
        RECT  42.9 164.4 43.8 165.3 ;
        RECT  45.9 164.4 46.8 165.3 ;
        RECT  42.9 164.85 43.8 172.35 ;
        RECT  43.35 164.4 46.35 165.3 ;
        RECT  45.9 162.15 46.8 164.85 ;
        RECT  47.7 177.9 48.9 179.1 ;
        RECT  44.7 174.6 45.9 175.8 ;
        RECT  39.0 170.25 51.0 171.15 ;
        RECT  39.0 155.55 51.0 156.45 ;
        RECT  41.1 156.0 42.0 158.85 ;
        RECT  41.1 168.3 42.0 170.7 ;
        RECT  48.15 156.0 49.05 158.85 ;
        RECT  43.35 156.0 44.25 158.85 ;
        RECT  48.15 167.85 49.05 170.7 ;
        RECT  48.9 161.1 51.0 162.0 ;
        RECT  45.9 164.4 51.0 165.3 ;
        RECT  39.0 163.5 43.35 164.4 ;
        RECT  48.0 166.65 49.2 167.85 ;
        RECT  45.6 166.65 46.8 167.85 ;
        RECT  45.6 166.65 46.8 167.85 ;
        RECT  43.2 166.65 44.4 167.85 ;
        RECT  48.0 157.65 49.2 158.85 ;
        RECT  45.6 157.65 46.8 158.85 ;
        RECT  45.6 157.65 46.8 158.85 ;
        RECT  43.2 157.65 44.4 158.85 ;
        RECT  40.8 157.65 42.0 158.85 ;
        RECT  40.8 167.85 42.0 169.05 ;
        RECT  42.9 161.1 43.8 162.0 ;
        RECT  45.9 161.1 46.8 162.0 ;
        RECT  42.9 161.55 43.8 169.05 ;
        RECT  43.35 161.1 46.35 162.0 ;
        RECT  45.9 158.85 46.8 161.55 ;
        RECT  47.7 161.1 48.9 162.3 ;
        RECT  44.7 164.4 45.9 165.6 ;
        RECT  39.0 199.65 51.0 200.55 ;
        RECT  39.0 214.35 51.0 215.25 ;
        RECT  41.1 211.95 42.0 214.8 ;
        RECT  41.1 200.1 42.0 202.5 ;
        RECT  48.15 211.95 49.05 214.8 ;
        RECT  43.35 211.95 44.25 214.8 ;
        RECT  48.15 200.1 49.05 202.95 ;
        RECT  48.9 208.8 51.0 209.7 ;
        RECT  45.9 205.5 51.0 206.4 ;
        RECT  39.0 206.4 43.35 207.3 ;
        RECT  48.0 206.55 49.2 207.75 ;
        RECT  45.6 206.55 46.8 207.75 ;
        RECT  45.6 206.55 46.8 207.75 ;
        RECT  43.2 206.55 44.4 207.75 ;
        RECT  48.0 205.95 49.2 207.15 ;
        RECT  45.6 205.95 46.8 207.15 ;
        RECT  45.6 205.95 46.8 207.15 ;
        RECT  43.2 205.95 44.4 207.15 ;
        RECT  40.8 210.75 42.0 211.95 ;
        RECT  40.8 200.55 42.0 201.75 ;
        RECT  42.9 193.8 43.8 194.7 ;
        RECT  45.9 193.8 46.8 194.7 ;
        RECT  42.9 194.25 43.8 201.75 ;
        RECT  43.35 193.8 46.35 194.7 ;
        RECT  45.9 191.55 46.8 194.25 ;
        RECT  47.7 207.3 48.9 208.5 ;
        RECT  44.7 204.0 45.9 205.2 ;
        RECT  58.2 151.65 59.4 152.85 ;
        RECT  77.4 146.4 78.6 147.6 ;
        RECT  56.1 157.05 57.3 158.25 ;
        RECT  75.3 162.3 76.5 163.5 ;
        RECT  58.2 148.8 59.4 150.0 ;
        RECT  56.1 145.5 57.3 146.7 ;
        RECT  54.0 159.9 55.2 161.1 ;
        RECT  56.1 163.2 57.3 164.4 ;
        RECT  58.2 178.2 59.4 179.4 ;
        RECT  51.9 174.9 53.1 176.1 ;
        RECT  54.0 189.3 55.2 190.5 ;
        RECT  77.4 189.3 78.6 190.5 ;
        RECT  51.9 192.6 53.1 193.8 ;
        RECT  75.3 192.6 76.5 193.8 ;
        RECT  60.3 139.65 61.5 140.85 ;
        RECT  62.4 154.35 63.6 155.55 ;
        RECT  60.3 169.05 61.5 170.25 ;
        RECT  62.4 183.75 63.6 184.95 ;
        RECT  60.3 196.2 61.5 197.4 ;
        RECT  29.4 199.65 41.4 200.55 ;
        RECT  29.4 214.35 41.4 215.25 ;
        RECT  38.4 211.95 39.3 214.8 ;
        RECT  38.4 200.1 39.3 202.5 ;
        RECT  31.35 211.95 32.25 214.8 ;
        RECT  36.15 211.95 37.05 214.8 ;
        RECT  31.35 200.1 32.25 202.95 ;
        RECT  29.4 208.8 31.5 209.7 ;
        RECT  29.4 205.5 34.5 206.4 ;
        RECT  37.05 206.4 41.4 207.3 ;
        RECT  31.2 202.95 32.4 204.15 ;
        RECT  33.6 202.95 34.8 204.15 ;
        RECT  33.6 202.95 34.8 204.15 ;
        RECT  36.0 202.95 37.2 204.15 ;
        RECT  31.2 211.95 32.4 213.15 ;
        RECT  33.6 211.95 34.8 213.15 ;
        RECT  33.6 211.95 34.8 213.15 ;
        RECT  36.0 211.95 37.2 213.15 ;
        RECT  38.4 211.95 39.6 213.15 ;
        RECT  38.4 201.75 39.6 202.95 ;
        RECT  36.6 208.8 37.5 209.7 ;
        RECT  33.6 208.8 34.5 209.7 ;
        RECT  36.6 201.75 37.5 209.25 ;
        RECT  34.05 208.8 37.05 209.7 ;
        RECT  33.6 209.25 34.5 211.95 ;
        RECT  31.5 208.5 32.7 209.7 ;
        RECT  34.5 205.2 35.7 206.4 ;
        RECT  29.4 229.05 41.4 229.95 ;
        RECT  29.4 214.35 41.4 215.25 ;
        RECT  38.4 214.8 39.3 217.65 ;
        RECT  38.4 227.1 39.3 229.5 ;
        RECT  31.35 214.8 32.25 217.65 ;
        RECT  36.15 214.8 37.05 217.65 ;
        RECT  31.35 226.65 32.25 229.5 ;
        RECT  29.4 219.9 31.5 220.8 ;
        RECT  29.4 223.2 34.5 224.1 ;
        RECT  37.05 222.3 41.4 223.2 ;
        RECT  31.2 221.85 32.4 223.05 ;
        RECT  33.6 221.85 34.8 223.05 ;
        RECT  33.6 221.85 34.8 223.05 ;
        RECT  36.0 221.85 37.2 223.05 ;
        RECT  31.2 222.45 32.4 223.65 ;
        RECT  33.6 222.45 34.8 223.65 ;
        RECT  33.6 222.45 34.8 223.65 ;
        RECT  36.0 222.45 37.2 223.65 ;
        RECT  38.4 217.65 39.6 218.85 ;
        RECT  38.4 227.85 39.6 229.05 ;
        RECT  36.6 234.9 37.5 235.8 ;
        RECT  33.6 234.9 34.5 235.8 ;
        RECT  36.6 227.85 37.5 235.35 ;
        RECT  34.05 234.9 37.05 235.8 ;
        RECT  33.6 235.35 34.5 238.05 ;
        RECT  31.5 221.1 32.7 222.3 ;
        RECT  34.5 224.4 35.7 225.6 ;
        RECT  29.4 229.05 41.4 229.95 ;
        RECT  29.4 243.75 41.4 244.65 ;
        RECT  38.4 241.35 39.3 244.2 ;
        RECT  38.4 229.5 39.3 231.9 ;
        RECT  31.35 241.35 32.25 244.2 ;
        RECT  36.15 241.35 37.05 244.2 ;
        RECT  31.35 229.5 32.25 232.35 ;
        RECT  29.4 238.2 31.5 239.1 ;
        RECT  29.4 234.9 34.5 235.8 ;
        RECT  37.05 235.8 41.4 236.7 ;
        RECT  31.2 232.35 32.4 233.55 ;
        RECT  33.6 232.35 34.8 233.55 ;
        RECT  33.6 232.35 34.8 233.55 ;
        RECT  36.0 232.35 37.2 233.55 ;
        RECT  31.2 241.35 32.4 242.55 ;
        RECT  33.6 241.35 34.8 242.55 ;
        RECT  33.6 241.35 34.8 242.55 ;
        RECT  36.0 241.35 37.2 242.55 ;
        RECT  38.4 241.35 39.6 242.55 ;
        RECT  38.4 231.15 39.6 232.35 ;
        RECT  36.6 238.2 37.5 239.1 ;
        RECT  33.6 238.2 34.5 239.1 ;
        RECT  36.6 231.15 37.5 238.65 ;
        RECT  34.05 238.2 37.05 239.1 ;
        RECT  33.6 238.65 34.5 241.35 ;
        RECT  31.5 237.9 32.7 239.1 ;
        RECT  34.5 234.6 35.7 235.8 ;
        RECT  29.4 258.45 41.4 259.35 ;
        RECT  29.4 243.75 41.4 244.65 ;
        RECT  38.4 244.2 39.3 247.05 ;
        RECT  38.4 256.5 39.3 258.9 ;
        RECT  31.35 244.2 32.25 247.05 ;
        RECT  36.15 244.2 37.05 247.05 ;
        RECT  31.35 256.05 32.25 258.9 ;
        RECT  29.4 249.3 31.5 250.2 ;
        RECT  29.4 252.6 34.5 253.5 ;
        RECT  37.05 251.7 41.4 252.6 ;
        RECT  31.2 251.25 32.4 252.45 ;
        RECT  33.6 251.25 34.8 252.45 ;
        RECT  33.6 251.25 34.8 252.45 ;
        RECT  36.0 251.25 37.2 252.45 ;
        RECT  31.2 251.85 32.4 253.05 ;
        RECT  33.6 251.85 34.8 253.05 ;
        RECT  33.6 251.85 34.8 253.05 ;
        RECT  36.0 251.85 37.2 253.05 ;
        RECT  38.4 247.05 39.6 248.25 ;
        RECT  38.4 257.25 39.6 258.45 ;
        RECT  36.6 264.3 37.5 265.2 ;
        RECT  33.6 264.3 34.5 265.2 ;
        RECT  36.6 257.25 37.5 264.75 ;
        RECT  34.05 264.3 37.05 265.2 ;
        RECT  33.6 264.75 34.5 267.45 ;
        RECT  31.5 250.5 32.7 251.7 ;
        RECT  34.5 253.8 35.7 255.0 ;
        RECT  29.4 258.45 41.4 259.35 ;
        RECT  29.4 273.15 41.4 274.05 ;
        RECT  38.4 270.75 39.3 273.6 ;
        RECT  38.4 258.9 39.3 261.3 ;
        RECT  31.35 270.75 32.25 273.6 ;
        RECT  36.15 270.75 37.05 273.6 ;
        RECT  31.35 258.9 32.25 261.75 ;
        RECT  29.4 267.6 31.5 268.5 ;
        RECT  29.4 264.3 34.5 265.2 ;
        RECT  37.05 265.2 41.4 266.1 ;
        RECT  31.2 261.75 32.4 262.95 ;
        RECT  33.6 261.75 34.8 262.95 ;
        RECT  33.6 261.75 34.8 262.95 ;
        RECT  36.0 261.75 37.2 262.95 ;
        RECT  31.2 270.75 32.4 271.95 ;
        RECT  33.6 270.75 34.8 271.95 ;
        RECT  33.6 270.75 34.8 271.95 ;
        RECT  36.0 270.75 37.2 271.95 ;
        RECT  38.4 270.75 39.6 271.95 ;
        RECT  38.4 260.55 39.6 261.75 ;
        RECT  36.6 267.6 37.5 268.5 ;
        RECT  33.6 267.6 34.5 268.5 ;
        RECT  36.6 260.55 37.5 268.05 ;
        RECT  34.05 267.6 37.05 268.5 ;
        RECT  33.6 268.05 34.5 270.75 ;
        RECT  31.5 267.3 32.7 268.5 ;
        RECT  34.5 264.0 35.7 265.2 ;
        RECT  29.4 287.85 41.4 288.75 ;
        RECT  29.4 273.15 41.4 274.05 ;
        RECT  38.4 273.6 39.3 276.45 ;
        RECT  38.4 285.9 39.3 288.3 ;
        RECT  31.35 273.6 32.25 276.45 ;
        RECT  36.15 273.6 37.05 276.45 ;
        RECT  31.35 285.45 32.25 288.3 ;
        RECT  29.4 278.7 31.5 279.6 ;
        RECT  29.4 282.0 34.5 282.9 ;
        RECT  37.05 281.1 41.4 282.0 ;
        RECT  31.2 280.65 32.4 281.85 ;
        RECT  33.6 280.65 34.8 281.85 ;
        RECT  33.6 280.65 34.8 281.85 ;
        RECT  36.0 280.65 37.2 281.85 ;
        RECT  31.2 281.25 32.4 282.45 ;
        RECT  33.6 281.25 34.8 282.45 ;
        RECT  33.6 281.25 34.8 282.45 ;
        RECT  36.0 281.25 37.2 282.45 ;
        RECT  38.4 276.45 39.6 277.65 ;
        RECT  38.4 286.65 39.6 287.85 ;
        RECT  36.6 293.7 37.5 294.6 ;
        RECT  33.6 293.7 34.5 294.6 ;
        RECT  36.6 286.65 37.5 294.15 ;
        RECT  34.05 293.7 37.05 294.6 ;
        RECT  33.6 294.15 34.5 296.85 ;
        RECT  31.5 279.9 32.7 281.1 ;
        RECT  34.5 283.2 35.7 284.4 ;
        RECT  29.4 287.85 41.4 288.75 ;
        RECT  29.4 302.55 41.4 303.45 ;
        RECT  38.4 300.15 39.3 303.0 ;
        RECT  38.4 288.3 39.3 290.7 ;
        RECT  31.35 300.15 32.25 303.0 ;
        RECT  36.15 300.15 37.05 303.0 ;
        RECT  31.35 288.3 32.25 291.15 ;
        RECT  29.4 297.0 31.5 297.9 ;
        RECT  29.4 293.7 34.5 294.6 ;
        RECT  37.05 294.6 41.4 295.5 ;
        RECT  31.2 291.15 32.4 292.35 ;
        RECT  33.6 291.15 34.8 292.35 ;
        RECT  33.6 291.15 34.8 292.35 ;
        RECT  36.0 291.15 37.2 292.35 ;
        RECT  31.2 300.15 32.4 301.35 ;
        RECT  33.6 300.15 34.8 301.35 ;
        RECT  33.6 300.15 34.8 301.35 ;
        RECT  36.0 300.15 37.2 301.35 ;
        RECT  38.4 300.15 39.6 301.35 ;
        RECT  38.4 289.95 39.6 291.15 ;
        RECT  36.6 297.0 37.5 297.9 ;
        RECT  33.6 297.0 34.5 297.9 ;
        RECT  36.6 289.95 37.5 297.45 ;
        RECT  34.05 297.0 37.05 297.9 ;
        RECT  33.6 297.45 34.5 300.15 ;
        RECT  31.5 296.7 32.7 297.9 ;
        RECT  34.5 293.4 35.7 294.6 ;
        RECT  29.4 317.25 41.4 318.15 ;
        RECT  29.4 302.55 41.4 303.45 ;
        RECT  38.4 303.0 39.3 305.85 ;
        RECT  38.4 315.3 39.3 317.7 ;
        RECT  31.35 303.0 32.25 305.85 ;
        RECT  36.15 303.0 37.05 305.85 ;
        RECT  31.35 314.85 32.25 317.7 ;
        RECT  29.4 308.1 31.5 309.0 ;
        RECT  29.4 311.4 34.5 312.3 ;
        RECT  37.05 310.5 41.4 311.4 ;
        RECT  31.2 310.05 32.4 311.25 ;
        RECT  33.6 310.05 34.8 311.25 ;
        RECT  33.6 310.05 34.8 311.25 ;
        RECT  36.0 310.05 37.2 311.25 ;
        RECT  31.2 310.65 32.4 311.85 ;
        RECT  33.6 310.65 34.8 311.85 ;
        RECT  33.6 310.65 34.8 311.85 ;
        RECT  36.0 310.65 37.2 311.85 ;
        RECT  38.4 305.85 39.6 307.05 ;
        RECT  38.4 316.05 39.6 317.25 ;
        RECT  36.6 323.1 37.5 324.0 ;
        RECT  33.6 323.1 34.5 324.0 ;
        RECT  36.6 316.05 37.5 323.55 ;
        RECT  34.05 323.1 37.05 324.0 ;
        RECT  33.6 323.55 34.5 326.25 ;
        RECT  31.5 309.3 32.7 310.5 ;
        RECT  34.5 312.6 35.7 313.8 ;
        RECT  29.4 317.25 41.4 318.15 ;
        RECT  29.4 331.95 41.4 332.85 ;
        RECT  38.4 329.55 39.3 332.4 ;
        RECT  38.4 317.7 39.3 320.1 ;
        RECT  31.35 329.55 32.25 332.4 ;
        RECT  36.15 329.55 37.05 332.4 ;
        RECT  31.35 317.7 32.25 320.55 ;
        RECT  29.4 326.4 31.5 327.3 ;
        RECT  29.4 323.1 34.5 324.0 ;
        RECT  37.05 324.0 41.4 324.9 ;
        RECT  31.2 320.55 32.4 321.75 ;
        RECT  33.6 320.55 34.8 321.75 ;
        RECT  33.6 320.55 34.8 321.75 ;
        RECT  36.0 320.55 37.2 321.75 ;
        RECT  31.2 329.55 32.4 330.75 ;
        RECT  33.6 329.55 34.8 330.75 ;
        RECT  33.6 329.55 34.8 330.75 ;
        RECT  36.0 329.55 37.2 330.75 ;
        RECT  38.4 329.55 39.6 330.75 ;
        RECT  38.4 319.35 39.6 320.55 ;
        RECT  36.6 326.4 37.5 327.3 ;
        RECT  33.6 326.4 34.5 327.3 ;
        RECT  36.6 319.35 37.5 326.85 ;
        RECT  34.05 326.4 37.05 327.3 ;
        RECT  33.6 326.85 34.5 329.55 ;
        RECT  31.5 326.1 32.7 327.3 ;
        RECT  34.5 322.8 35.7 324.0 ;
        RECT  29.4 346.65 41.4 347.55 ;
        RECT  29.4 331.95 41.4 332.85 ;
        RECT  38.4 332.4 39.3 335.25 ;
        RECT  38.4 344.7 39.3 347.1 ;
        RECT  31.35 332.4 32.25 335.25 ;
        RECT  36.15 332.4 37.05 335.25 ;
        RECT  31.35 344.25 32.25 347.1 ;
        RECT  29.4 337.5 31.5 338.4 ;
        RECT  29.4 340.8 34.5 341.7 ;
        RECT  37.05 339.9 41.4 340.8 ;
        RECT  31.2 339.45 32.4 340.65 ;
        RECT  33.6 339.45 34.8 340.65 ;
        RECT  33.6 339.45 34.8 340.65 ;
        RECT  36.0 339.45 37.2 340.65 ;
        RECT  31.2 340.05 32.4 341.25 ;
        RECT  33.6 340.05 34.8 341.25 ;
        RECT  33.6 340.05 34.8 341.25 ;
        RECT  36.0 340.05 37.2 341.25 ;
        RECT  38.4 335.25 39.6 336.45 ;
        RECT  38.4 345.45 39.6 346.65 ;
        RECT  36.6 352.5 37.5 353.4 ;
        RECT  33.6 352.5 34.5 353.4 ;
        RECT  36.6 345.45 37.5 352.95 ;
        RECT  34.05 352.5 37.05 353.4 ;
        RECT  33.6 352.95 34.5 355.65 ;
        RECT  31.5 338.7 32.7 339.9 ;
        RECT  34.5 342.0 35.7 343.2 ;
        RECT  29.4 346.65 41.4 347.55 ;
        RECT  29.4 361.35 41.4 362.25 ;
        RECT  38.4 358.95 39.3 361.8 ;
        RECT  38.4 347.1 39.3 349.5 ;
        RECT  31.35 358.95 32.25 361.8 ;
        RECT  36.15 358.95 37.05 361.8 ;
        RECT  31.35 347.1 32.25 349.95 ;
        RECT  29.4 355.8 31.5 356.7 ;
        RECT  29.4 352.5 34.5 353.4 ;
        RECT  37.05 353.4 41.4 354.3 ;
        RECT  31.2 349.95 32.4 351.15 ;
        RECT  33.6 349.95 34.8 351.15 ;
        RECT  33.6 349.95 34.8 351.15 ;
        RECT  36.0 349.95 37.2 351.15 ;
        RECT  31.2 358.95 32.4 360.15 ;
        RECT  33.6 358.95 34.8 360.15 ;
        RECT  33.6 358.95 34.8 360.15 ;
        RECT  36.0 358.95 37.2 360.15 ;
        RECT  38.4 358.95 39.6 360.15 ;
        RECT  38.4 348.75 39.6 349.95 ;
        RECT  36.6 355.8 37.5 356.7 ;
        RECT  33.6 355.8 34.5 356.7 ;
        RECT  36.6 348.75 37.5 356.25 ;
        RECT  34.05 355.8 37.05 356.7 ;
        RECT  33.6 356.25 34.5 358.95 ;
        RECT  31.5 355.5 32.7 356.7 ;
        RECT  34.5 352.2 35.7 353.4 ;
        RECT  29.4 376.05 41.4 376.95 ;
        RECT  29.4 361.35 41.4 362.25 ;
        RECT  38.4 361.8 39.3 364.65 ;
        RECT  38.4 374.1 39.3 376.5 ;
        RECT  31.35 361.8 32.25 364.65 ;
        RECT  36.15 361.8 37.05 364.65 ;
        RECT  31.35 373.65 32.25 376.5 ;
        RECT  29.4 366.9 31.5 367.8 ;
        RECT  29.4 370.2 34.5 371.1 ;
        RECT  37.05 369.3 41.4 370.2 ;
        RECT  31.2 368.85 32.4 370.05 ;
        RECT  33.6 368.85 34.8 370.05 ;
        RECT  33.6 368.85 34.8 370.05 ;
        RECT  36.0 368.85 37.2 370.05 ;
        RECT  31.2 369.45 32.4 370.65 ;
        RECT  33.6 369.45 34.8 370.65 ;
        RECT  33.6 369.45 34.8 370.65 ;
        RECT  36.0 369.45 37.2 370.65 ;
        RECT  38.4 364.65 39.6 365.85 ;
        RECT  38.4 374.85 39.6 376.05 ;
        RECT  36.6 381.9 37.5 382.8 ;
        RECT  33.6 381.9 34.5 382.8 ;
        RECT  36.6 374.85 37.5 382.35 ;
        RECT  34.05 381.9 37.05 382.8 ;
        RECT  33.6 382.35 34.5 385.05 ;
        RECT  31.5 368.1 32.7 369.3 ;
        RECT  34.5 371.4 35.7 372.6 ;
        RECT  29.4 376.05 41.4 376.95 ;
        RECT  29.4 390.75 41.4 391.65 ;
        RECT  38.4 388.35 39.3 391.2 ;
        RECT  38.4 376.5 39.3 378.9 ;
        RECT  31.35 388.35 32.25 391.2 ;
        RECT  36.15 388.35 37.05 391.2 ;
        RECT  31.35 376.5 32.25 379.35 ;
        RECT  29.4 385.2 31.5 386.1 ;
        RECT  29.4 381.9 34.5 382.8 ;
        RECT  37.05 382.8 41.4 383.7 ;
        RECT  31.2 379.35 32.4 380.55 ;
        RECT  33.6 379.35 34.8 380.55 ;
        RECT  33.6 379.35 34.8 380.55 ;
        RECT  36.0 379.35 37.2 380.55 ;
        RECT  31.2 388.35 32.4 389.55 ;
        RECT  33.6 388.35 34.8 389.55 ;
        RECT  33.6 388.35 34.8 389.55 ;
        RECT  36.0 388.35 37.2 389.55 ;
        RECT  38.4 388.35 39.6 389.55 ;
        RECT  38.4 378.15 39.6 379.35 ;
        RECT  36.6 385.2 37.5 386.1 ;
        RECT  33.6 385.2 34.5 386.1 ;
        RECT  36.6 378.15 37.5 385.65 ;
        RECT  34.05 385.2 37.05 386.1 ;
        RECT  33.6 385.65 34.5 388.35 ;
        RECT  31.5 384.9 32.7 386.1 ;
        RECT  34.5 381.6 35.7 382.8 ;
        RECT  29.4 405.45 41.4 406.35 ;
        RECT  29.4 390.75 41.4 391.65 ;
        RECT  38.4 391.2 39.3 394.05 ;
        RECT  38.4 403.5 39.3 405.9 ;
        RECT  31.35 391.2 32.25 394.05 ;
        RECT  36.15 391.2 37.05 394.05 ;
        RECT  31.35 403.05 32.25 405.9 ;
        RECT  29.4 396.3 31.5 397.2 ;
        RECT  29.4 399.6 34.5 400.5 ;
        RECT  37.05 398.7 41.4 399.6 ;
        RECT  31.2 398.25 32.4 399.45 ;
        RECT  33.6 398.25 34.8 399.45 ;
        RECT  33.6 398.25 34.8 399.45 ;
        RECT  36.0 398.25 37.2 399.45 ;
        RECT  31.2 398.85 32.4 400.05 ;
        RECT  33.6 398.85 34.8 400.05 ;
        RECT  33.6 398.85 34.8 400.05 ;
        RECT  36.0 398.85 37.2 400.05 ;
        RECT  38.4 394.05 39.6 395.25 ;
        RECT  38.4 404.25 39.6 405.45 ;
        RECT  36.6 411.3 37.5 412.2 ;
        RECT  33.6 411.3 34.5 412.2 ;
        RECT  36.6 404.25 37.5 411.75 ;
        RECT  34.05 411.3 37.05 412.2 ;
        RECT  33.6 411.75 34.5 414.45 ;
        RECT  31.5 397.5 32.7 398.7 ;
        RECT  34.5 400.8 35.7 402.0 ;
        RECT  29.4 405.45 41.4 406.35 ;
        RECT  29.4 420.15 41.4 421.05 ;
        RECT  38.4 417.75 39.3 420.6 ;
        RECT  38.4 405.9 39.3 408.3 ;
        RECT  31.35 417.75 32.25 420.6 ;
        RECT  36.15 417.75 37.05 420.6 ;
        RECT  31.35 405.9 32.25 408.75 ;
        RECT  29.4 414.6 31.5 415.5 ;
        RECT  29.4 411.3 34.5 412.2 ;
        RECT  37.05 412.2 41.4 413.1 ;
        RECT  31.2 408.75 32.4 409.95 ;
        RECT  33.6 408.75 34.8 409.95 ;
        RECT  33.6 408.75 34.8 409.95 ;
        RECT  36.0 408.75 37.2 409.95 ;
        RECT  31.2 417.75 32.4 418.95 ;
        RECT  33.6 417.75 34.8 418.95 ;
        RECT  33.6 417.75 34.8 418.95 ;
        RECT  36.0 417.75 37.2 418.95 ;
        RECT  38.4 417.75 39.6 418.95 ;
        RECT  38.4 407.55 39.6 408.75 ;
        RECT  36.6 414.6 37.5 415.5 ;
        RECT  33.6 414.6 34.5 415.5 ;
        RECT  36.6 407.55 37.5 415.05 ;
        RECT  34.05 414.6 37.05 415.5 ;
        RECT  33.6 415.05 34.5 417.75 ;
        RECT  31.5 414.3 32.7 415.5 ;
        RECT  34.5 411.0 35.7 412.2 ;
        RECT  29.4 434.85 41.4 435.75 ;
        RECT  29.4 420.15 41.4 421.05 ;
        RECT  38.4 420.6 39.3 423.45 ;
        RECT  38.4 432.9 39.3 435.3 ;
        RECT  31.35 420.6 32.25 423.45 ;
        RECT  36.15 420.6 37.05 423.45 ;
        RECT  31.35 432.45 32.25 435.3 ;
        RECT  29.4 425.7 31.5 426.6 ;
        RECT  29.4 429.0 34.5 429.9 ;
        RECT  37.05 428.1 41.4 429.0 ;
        RECT  31.2 427.65 32.4 428.85 ;
        RECT  33.6 427.65 34.8 428.85 ;
        RECT  33.6 427.65 34.8 428.85 ;
        RECT  36.0 427.65 37.2 428.85 ;
        RECT  31.2 428.25 32.4 429.45 ;
        RECT  33.6 428.25 34.8 429.45 ;
        RECT  33.6 428.25 34.8 429.45 ;
        RECT  36.0 428.25 37.2 429.45 ;
        RECT  38.4 423.45 39.6 424.65 ;
        RECT  38.4 433.65 39.6 434.85 ;
        RECT  36.6 440.7 37.5 441.6 ;
        RECT  33.6 440.7 34.5 441.6 ;
        RECT  36.6 433.65 37.5 441.15 ;
        RECT  34.05 440.7 37.05 441.6 ;
        RECT  33.6 441.15 34.5 443.85 ;
        RECT  31.5 426.9 32.7 428.1 ;
        RECT  34.5 430.2 35.7 431.4 ;
        RECT  41.4 199.65 51.0 200.55 ;
        RECT  41.4 214.35 51.0 215.25 ;
        RECT  48.0 211.95 49.2 214.35 ;
        RECT  48.0 200.55 49.2 202.35 ;
        RECT  43.2 200.55 44.4 201.45 ;
        RECT  43.2 213.15 44.4 214.35 ;
        RECT  45.6 202.65 46.8 212.1 ;
        RECT  41.4 206.4 43.5 207.3 ;
        RECT  46.8 206.4 51.0 207.3 ;
        RECT  43.2 202.65 44.4 203.85 ;
        RECT  45.6 202.65 46.8 203.85 ;
        RECT  43.2 211.95 44.4 213.15 ;
        RECT  45.6 211.95 46.8 213.15 ;
        RECT  48.0 211.95 49.2 213.15 ;
        RECT  48.0 201.45 49.2 202.65 ;
        RECT  43.5 206.25 44.7 207.45 ;
        RECT  41.4 229.05 51.0 229.95 ;
        RECT  41.4 214.35 51.0 215.25 ;
        RECT  48.0 215.25 49.2 217.65 ;
        RECT  48.0 227.25 49.2 229.05 ;
        RECT  43.2 228.15 44.4 229.05 ;
        RECT  43.2 215.25 44.4 216.45 ;
        RECT  45.6 217.5 46.8 226.95 ;
        RECT  41.4 222.3 43.5 223.2 ;
        RECT  46.8 222.3 51.0 223.2 ;
        RECT  43.2 223.35 44.4 224.55 ;
        RECT  45.6 223.35 46.8 224.55 ;
        RECT  43.2 222.45 44.4 223.65 ;
        RECT  45.6 222.45 46.8 223.65 ;
        RECT  48.0 217.65 49.2 218.85 ;
        RECT  48.0 228.15 49.2 229.35 ;
        RECT  43.5 223.35 44.7 224.55 ;
        RECT  41.4 229.05 51.0 229.95 ;
        RECT  41.4 243.75 51.0 244.65 ;
        RECT  48.0 241.35 49.2 243.75 ;
        RECT  48.0 229.95 49.2 231.75 ;
        RECT  43.2 229.95 44.4 230.85 ;
        RECT  43.2 242.55 44.4 243.75 ;
        RECT  45.6 232.05 46.8 241.5 ;
        RECT  41.4 235.8 43.5 236.7 ;
        RECT  46.8 235.8 51.0 236.7 ;
        RECT  43.2 232.05 44.4 233.25 ;
        RECT  45.6 232.05 46.8 233.25 ;
        RECT  43.2 241.35 44.4 242.55 ;
        RECT  45.6 241.35 46.8 242.55 ;
        RECT  48.0 241.35 49.2 242.55 ;
        RECT  48.0 230.85 49.2 232.05 ;
        RECT  43.5 235.65 44.7 236.85 ;
        RECT  41.4 258.45 51.0 259.35 ;
        RECT  41.4 243.75 51.0 244.65 ;
        RECT  48.0 244.65 49.2 247.05 ;
        RECT  48.0 256.65 49.2 258.45 ;
        RECT  43.2 257.55 44.4 258.45 ;
        RECT  43.2 244.65 44.4 245.85 ;
        RECT  45.6 246.9 46.8 256.35 ;
        RECT  41.4 251.7 43.5 252.6 ;
        RECT  46.8 251.7 51.0 252.6 ;
        RECT  43.2 252.75 44.4 253.95 ;
        RECT  45.6 252.75 46.8 253.95 ;
        RECT  43.2 251.85 44.4 253.05 ;
        RECT  45.6 251.85 46.8 253.05 ;
        RECT  48.0 247.05 49.2 248.25 ;
        RECT  48.0 257.55 49.2 258.75 ;
        RECT  43.5 252.75 44.7 253.95 ;
        RECT  41.4 258.45 51.0 259.35 ;
        RECT  41.4 273.15 51.0 274.05 ;
        RECT  48.0 270.75 49.2 273.15 ;
        RECT  48.0 259.35 49.2 261.15 ;
        RECT  43.2 259.35 44.4 260.25 ;
        RECT  43.2 271.95 44.4 273.15 ;
        RECT  45.6 261.45 46.8 270.9 ;
        RECT  41.4 265.2 43.5 266.1 ;
        RECT  46.8 265.2 51.0 266.1 ;
        RECT  43.2 261.45 44.4 262.65 ;
        RECT  45.6 261.45 46.8 262.65 ;
        RECT  43.2 270.75 44.4 271.95 ;
        RECT  45.6 270.75 46.8 271.95 ;
        RECT  48.0 270.75 49.2 271.95 ;
        RECT  48.0 260.25 49.2 261.45 ;
        RECT  43.5 265.05 44.7 266.25 ;
        RECT  41.4 287.85 51.0 288.75 ;
        RECT  41.4 273.15 51.0 274.05 ;
        RECT  48.0 274.05 49.2 276.45 ;
        RECT  48.0 286.05 49.2 287.85 ;
        RECT  43.2 286.95 44.4 287.85 ;
        RECT  43.2 274.05 44.4 275.25 ;
        RECT  45.6 276.3 46.8 285.75 ;
        RECT  41.4 281.1 43.5 282.0 ;
        RECT  46.8 281.1 51.0 282.0 ;
        RECT  43.2 282.15 44.4 283.35 ;
        RECT  45.6 282.15 46.8 283.35 ;
        RECT  43.2 281.25 44.4 282.45 ;
        RECT  45.6 281.25 46.8 282.45 ;
        RECT  48.0 276.45 49.2 277.65 ;
        RECT  48.0 286.95 49.2 288.15 ;
        RECT  43.5 282.15 44.7 283.35 ;
        RECT  41.4 287.85 51.0 288.75 ;
        RECT  41.4 302.55 51.0 303.45 ;
        RECT  48.0 300.15 49.2 302.55 ;
        RECT  48.0 288.75 49.2 290.55 ;
        RECT  43.2 288.75 44.4 289.65 ;
        RECT  43.2 301.35 44.4 302.55 ;
        RECT  45.6 290.85 46.8 300.3 ;
        RECT  41.4 294.6 43.5 295.5 ;
        RECT  46.8 294.6 51.0 295.5 ;
        RECT  43.2 290.85 44.4 292.05 ;
        RECT  45.6 290.85 46.8 292.05 ;
        RECT  43.2 300.15 44.4 301.35 ;
        RECT  45.6 300.15 46.8 301.35 ;
        RECT  48.0 300.15 49.2 301.35 ;
        RECT  48.0 289.65 49.2 290.85 ;
        RECT  43.5 294.45 44.7 295.65 ;
        RECT  41.4 317.25 51.0 318.15 ;
        RECT  41.4 302.55 51.0 303.45 ;
        RECT  48.0 303.45 49.2 305.85 ;
        RECT  48.0 315.45 49.2 317.25 ;
        RECT  43.2 316.35 44.4 317.25 ;
        RECT  43.2 303.45 44.4 304.65 ;
        RECT  45.6 305.7 46.8 315.15 ;
        RECT  41.4 310.5 43.5 311.4 ;
        RECT  46.8 310.5 51.0 311.4 ;
        RECT  43.2 311.55 44.4 312.75 ;
        RECT  45.6 311.55 46.8 312.75 ;
        RECT  43.2 310.65 44.4 311.85 ;
        RECT  45.6 310.65 46.8 311.85 ;
        RECT  48.0 305.85 49.2 307.05 ;
        RECT  48.0 316.35 49.2 317.55 ;
        RECT  43.5 311.55 44.7 312.75 ;
        RECT  41.4 317.25 51.0 318.15 ;
        RECT  41.4 331.95 51.0 332.85 ;
        RECT  48.0 329.55 49.2 331.95 ;
        RECT  48.0 318.15 49.2 319.95 ;
        RECT  43.2 318.15 44.4 319.05 ;
        RECT  43.2 330.75 44.4 331.95 ;
        RECT  45.6 320.25 46.8 329.7 ;
        RECT  41.4 324.0 43.5 324.9 ;
        RECT  46.8 324.0 51.0 324.9 ;
        RECT  43.2 320.25 44.4 321.45 ;
        RECT  45.6 320.25 46.8 321.45 ;
        RECT  43.2 329.55 44.4 330.75 ;
        RECT  45.6 329.55 46.8 330.75 ;
        RECT  48.0 329.55 49.2 330.75 ;
        RECT  48.0 319.05 49.2 320.25 ;
        RECT  43.5 323.85 44.7 325.05 ;
        RECT  41.4 346.65 51.0 347.55 ;
        RECT  41.4 331.95 51.0 332.85 ;
        RECT  48.0 332.85 49.2 335.25 ;
        RECT  48.0 344.85 49.2 346.65 ;
        RECT  43.2 345.75 44.4 346.65 ;
        RECT  43.2 332.85 44.4 334.05 ;
        RECT  45.6 335.1 46.8 344.55 ;
        RECT  41.4 339.9 43.5 340.8 ;
        RECT  46.8 339.9 51.0 340.8 ;
        RECT  43.2 340.95 44.4 342.15 ;
        RECT  45.6 340.95 46.8 342.15 ;
        RECT  43.2 340.05 44.4 341.25 ;
        RECT  45.6 340.05 46.8 341.25 ;
        RECT  48.0 335.25 49.2 336.45 ;
        RECT  48.0 345.75 49.2 346.95 ;
        RECT  43.5 340.95 44.7 342.15 ;
        RECT  41.4 346.65 51.0 347.55 ;
        RECT  41.4 361.35 51.0 362.25 ;
        RECT  48.0 358.95 49.2 361.35 ;
        RECT  48.0 347.55 49.2 349.35 ;
        RECT  43.2 347.55 44.4 348.45 ;
        RECT  43.2 360.15 44.4 361.35 ;
        RECT  45.6 349.65 46.8 359.1 ;
        RECT  41.4 353.4 43.5 354.3 ;
        RECT  46.8 353.4 51.0 354.3 ;
        RECT  43.2 349.65 44.4 350.85 ;
        RECT  45.6 349.65 46.8 350.85 ;
        RECT  43.2 358.95 44.4 360.15 ;
        RECT  45.6 358.95 46.8 360.15 ;
        RECT  48.0 358.95 49.2 360.15 ;
        RECT  48.0 348.45 49.2 349.65 ;
        RECT  43.5 353.25 44.7 354.45 ;
        RECT  41.4 376.05 51.0 376.95 ;
        RECT  41.4 361.35 51.0 362.25 ;
        RECT  48.0 362.25 49.2 364.65 ;
        RECT  48.0 374.25 49.2 376.05 ;
        RECT  43.2 375.15 44.4 376.05 ;
        RECT  43.2 362.25 44.4 363.45 ;
        RECT  45.6 364.5 46.8 373.95 ;
        RECT  41.4 369.3 43.5 370.2 ;
        RECT  46.8 369.3 51.0 370.2 ;
        RECT  43.2 370.35 44.4 371.55 ;
        RECT  45.6 370.35 46.8 371.55 ;
        RECT  43.2 369.45 44.4 370.65 ;
        RECT  45.6 369.45 46.8 370.65 ;
        RECT  48.0 364.65 49.2 365.85 ;
        RECT  48.0 375.15 49.2 376.35 ;
        RECT  43.5 370.35 44.7 371.55 ;
        RECT  41.4 376.05 51.0 376.95 ;
        RECT  41.4 390.75 51.0 391.65 ;
        RECT  48.0 388.35 49.2 390.75 ;
        RECT  48.0 376.95 49.2 378.75 ;
        RECT  43.2 376.95 44.4 377.85 ;
        RECT  43.2 389.55 44.4 390.75 ;
        RECT  45.6 379.05 46.8 388.5 ;
        RECT  41.4 382.8 43.5 383.7 ;
        RECT  46.8 382.8 51.0 383.7 ;
        RECT  43.2 379.05 44.4 380.25 ;
        RECT  45.6 379.05 46.8 380.25 ;
        RECT  43.2 388.35 44.4 389.55 ;
        RECT  45.6 388.35 46.8 389.55 ;
        RECT  48.0 388.35 49.2 389.55 ;
        RECT  48.0 377.85 49.2 379.05 ;
        RECT  43.5 382.65 44.7 383.85 ;
        RECT  41.4 405.45 51.0 406.35 ;
        RECT  41.4 390.75 51.0 391.65 ;
        RECT  48.0 391.65 49.2 394.05 ;
        RECT  48.0 403.65 49.2 405.45 ;
        RECT  43.2 404.55 44.4 405.45 ;
        RECT  43.2 391.65 44.4 392.85 ;
        RECT  45.6 393.9 46.8 403.35 ;
        RECT  41.4 398.7 43.5 399.6 ;
        RECT  46.8 398.7 51.0 399.6 ;
        RECT  43.2 399.75 44.4 400.95 ;
        RECT  45.6 399.75 46.8 400.95 ;
        RECT  43.2 398.85 44.4 400.05 ;
        RECT  45.6 398.85 46.8 400.05 ;
        RECT  48.0 394.05 49.2 395.25 ;
        RECT  48.0 404.55 49.2 405.75 ;
        RECT  43.5 399.75 44.7 400.95 ;
        RECT  41.4 405.45 51.0 406.35 ;
        RECT  41.4 420.15 51.0 421.05 ;
        RECT  48.0 417.75 49.2 420.15 ;
        RECT  48.0 406.35 49.2 408.15 ;
        RECT  43.2 406.35 44.4 407.25 ;
        RECT  43.2 418.95 44.4 420.15 ;
        RECT  45.6 408.45 46.8 417.9 ;
        RECT  41.4 412.2 43.5 413.1 ;
        RECT  46.8 412.2 51.0 413.1 ;
        RECT  43.2 408.45 44.4 409.65 ;
        RECT  45.6 408.45 46.8 409.65 ;
        RECT  43.2 417.75 44.4 418.95 ;
        RECT  45.6 417.75 46.8 418.95 ;
        RECT  48.0 417.75 49.2 418.95 ;
        RECT  48.0 407.25 49.2 408.45 ;
        RECT  43.5 412.05 44.7 413.25 ;
        RECT  41.4 434.85 51.0 435.75 ;
        RECT  41.4 420.15 51.0 421.05 ;
        RECT  48.0 421.05 49.2 423.45 ;
        RECT  48.0 433.05 49.2 434.85 ;
        RECT  43.2 433.95 44.4 434.85 ;
        RECT  43.2 421.05 44.4 422.25 ;
        RECT  45.6 423.3 46.8 432.75 ;
        RECT  41.4 428.1 43.5 429.0 ;
        RECT  46.8 428.1 51.0 429.0 ;
        RECT  43.2 429.15 44.4 430.35 ;
        RECT  45.6 429.15 46.8 430.35 ;
        RECT  43.2 428.25 44.4 429.45 ;
        RECT  45.6 428.25 46.8 429.45 ;
        RECT  48.0 423.45 49.2 424.65 ;
        RECT  48.0 433.95 49.2 435.15 ;
        RECT  43.5 429.15 44.7 430.35 ;
        RECT  12.6 88.8 13.8 90.0 ;
        RECT  14.7 104.7 15.9 105.9 ;
        RECT  16.8 118.2 18.0 119.4 ;
        RECT  18.9 134.1 20.1 135.3 ;
        RECT  21.0 147.6 22.2 148.8 ;
        RECT  23.1 163.5 24.3 164.7 ;
        RECT  25.2 177.0 26.4 178.2 ;
        RECT  27.3 192.9 28.5 194.1 ;
        RECT  12.6 208.8 13.8 210.0 ;
        RECT  21.0 205.5 22.2 206.7 ;
        RECT  12.6 219.9 13.8 221.1 ;
        RECT  23.1 223.2 24.3 224.4 ;
        RECT  12.6 238.2 13.8 239.4 ;
        RECT  25.2 234.9 26.4 236.1 ;
        RECT  12.6 249.3 13.8 250.5 ;
        RECT  27.3 252.6 28.5 253.8 ;
        RECT  14.7 267.6 15.9 268.8 ;
        RECT  21.0 264.3 22.2 265.5 ;
        RECT  14.7 278.7 15.9 279.9 ;
        RECT  23.1 282.0 24.3 283.2 ;
        RECT  14.7 297.0 15.9 298.2 ;
        RECT  25.2 293.7 26.4 294.9 ;
        RECT  14.7 308.1 15.9 309.3 ;
        RECT  27.3 311.4 28.5 312.6 ;
        RECT  16.8 326.4 18.0 327.6 ;
        RECT  21.0 323.1 22.2 324.3 ;
        RECT  16.8 337.5 18.0 338.7 ;
        RECT  23.1 340.8 24.3 342.0 ;
        RECT  16.8 355.8 18.0 357.0 ;
        RECT  25.2 352.5 26.4 353.7 ;
        RECT  16.8 366.9 18.0 368.1 ;
        RECT  27.3 370.2 28.5 371.4 ;
        RECT  18.9 385.2 20.1 386.4 ;
        RECT  21.0 381.9 22.2 383.1 ;
        RECT  18.9 396.3 20.1 397.5 ;
        RECT  23.1 399.6 24.3 400.8 ;
        RECT  18.9 414.6 20.1 415.8 ;
        RECT  25.2 411.3 26.4 412.5 ;
        RECT  18.9 425.7 20.1 426.9 ;
        RECT  27.3 429.0 28.5 430.2 ;
        RECT  53.7 201.9 54.6 440.7 ;
        RECT  53.7 206.4 58.2 207.3 ;
        RECT  66.0 205.5 66.9 207.3 ;
        RECT  78.9 206.4 79.8 207.3 ;
        RECT  88.5 206.4 89.4 207.3 ;
        RECT  53.7 222.3 58.2 223.2 ;
        RECT  66.0 222.3 66.9 224.1 ;
        RECT  78.9 222.3 79.8 223.2 ;
        RECT  87.6 222.3 88.5 223.2 ;
        RECT  53.7 235.8 58.2 236.7 ;
        RECT  66.0 234.9 66.9 236.7 ;
        RECT  78.9 235.8 79.8 236.7 ;
        RECT  88.5 235.8 89.4 236.7 ;
        RECT  53.7 251.7 58.2 252.6 ;
        RECT  66.0 251.7 66.9 253.5 ;
        RECT  78.9 251.7 79.8 252.6 ;
        RECT  87.6 251.7 88.5 252.6 ;
        RECT  53.7 265.2 58.2 266.1 ;
        RECT  66.0 264.3 66.9 266.1 ;
        RECT  78.9 265.2 79.8 266.1 ;
        RECT  88.5 265.2 89.4 266.1 ;
        RECT  53.7 281.1 58.2 282.0 ;
        RECT  66.0 281.1 66.9 282.9 ;
        RECT  78.9 281.1 79.8 282.0 ;
        RECT  87.6 281.1 88.5 282.0 ;
        RECT  53.7 294.6 58.2 295.5 ;
        RECT  66.0 293.7 66.9 295.5 ;
        RECT  78.9 294.6 79.8 295.5 ;
        RECT  88.5 294.6 89.4 295.5 ;
        RECT  53.7 310.5 58.2 311.4 ;
        RECT  66.0 310.5 66.9 312.3 ;
        RECT  78.9 310.5 79.8 311.4 ;
        RECT  87.6 310.5 88.5 311.4 ;
        RECT  53.7 324.0 58.2 324.9 ;
        RECT  66.0 323.1 66.9 324.9 ;
        RECT  78.9 324.0 79.8 324.9 ;
        RECT  88.5 324.0 89.4 324.9 ;
        RECT  53.7 339.9 58.2 340.8 ;
        RECT  66.0 339.9 66.9 341.7 ;
        RECT  78.9 339.9 79.8 340.8 ;
        RECT  87.6 339.9 88.5 340.8 ;
        RECT  53.7 353.4 58.2 354.3 ;
        RECT  66.0 352.5 66.9 354.3 ;
        RECT  78.9 353.4 79.8 354.3 ;
        RECT  88.5 353.4 89.4 354.3 ;
        RECT  53.7 369.3 58.2 370.2 ;
        RECT  66.0 369.3 66.9 371.1 ;
        RECT  78.9 369.3 79.8 370.2 ;
        RECT  87.6 369.3 88.5 370.2 ;
        RECT  53.7 382.8 58.2 383.7 ;
        RECT  66.0 381.9 66.9 383.7 ;
        RECT  78.9 382.8 79.8 383.7 ;
        RECT  88.5 382.8 89.4 383.7 ;
        RECT  53.7 398.7 58.2 399.6 ;
        RECT  66.0 398.7 66.9 400.5 ;
        RECT  78.9 398.7 79.8 399.6 ;
        RECT  87.6 398.7 88.5 399.6 ;
        RECT  53.7 412.2 58.2 413.1 ;
        RECT  66.0 411.3 66.9 413.1 ;
        RECT  78.9 412.2 79.8 413.1 ;
        RECT  88.5 412.2 89.4 413.1 ;
        RECT  53.7 428.1 58.2 429.0 ;
        RECT  66.0 428.1 66.9 429.9 ;
        RECT  78.9 428.1 79.8 429.0 ;
        RECT  87.6 428.1 88.5 429.0 ;
        RECT  50.7 214.35 51.9 215.55 ;
        RECT  57.0 214.35 58.2 215.55 ;
        RECT  57.3 199.65 66.9 200.55 ;
        RECT  57.3 214.35 66.9 215.25 ;
        RECT  63.9 211.95 65.1 214.35 ;
        RECT  63.9 200.55 65.1 202.35 ;
        RECT  59.1 200.55 60.3 201.45 ;
        RECT  59.1 213.15 60.3 214.35 ;
        RECT  61.5 202.65 62.7 212.1 ;
        RECT  57.3 206.4 59.4 207.3 ;
        RECT  62.7 206.4 66.9 207.3 ;
        RECT  59.1 202.65 60.3 203.85 ;
        RECT  61.5 202.65 62.7 203.85 ;
        RECT  59.1 211.95 60.3 213.15 ;
        RECT  61.5 211.95 62.7 213.15 ;
        RECT  63.9 211.95 65.1 213.15 ;
        RECT  63.9 201.45 65.1 202.65 ;
        RECT  59.4 206.25 60.6 207.45 ;
        RECT  66.9 199.65 78.9 200.55 ;
        RECT  66.9 214.35 78.9 215.25 ;
        RECT  75.9 211.95 76.8 214.8 ;
        RECT  75.9 200.1 76.8 202.5 ;
        RECT  68.85 211.95 69.75 214.8 ;
        RECT  73.65 211.95 74.55 214.8 ;
        RECT  68.85 200.1 69.75 202.95 ;
        RECT  66.9 208.8 69.0 209.7 ;
        RECT  66.9 205.5 72.0 206.4 ;
        RECT  74.55 206.4 78.9 207.3 ;
        RECT  68.7 202.95 69.9 204.15 ;
        RECT  71.1 202.95 72.3 204.15 ;
        RECT  71.1 202.95 72.3 204.15 ;
        RECT  73.5 202.95 74.7 204.15 ;
        RECT  68.7 211.95 69.9 213.15 ;
        RECT  71.1 211.95 72.3 213.15 ;
        RECT  71.1 211.95 72.3 213.15 ;
        RECT  73.5 211.95 74.7 213.15 ;
        RECT  75.9 211.95 77.1 213.15 ;
        RECT  75.9 201.75 77.1 202.95 ;
        RECT  74.1 208.8 75.0 209.7 ;
        RECT  71.1 208.8 72.0 209.7 ;
        RECT  74.1 201.75 75.0 209.25 ;
        RECT  71.55 208.8 74.55 209.7 ;
        RECT  71.1 209.25 72.0 211.95 ;
        RECT  69.0 208.5 70.2 209.7 ;
        RECT  72.0 205.2 73.2 206.4 ;
        RECT  78.9 199.65 88.5 200.55 ;
        RECT  78.9 214.35 88.5 215.25 ;
        RECT  85.5 211.95 86.7 214.35 ;
        RECT  85.5 200.55 86.7 202.35 ;
        RECT  80.7 200.55 81.9 201.45 ;
        RECT  80.7 213.15 81.9 214.35 ;
        RECT  83.1 202.65 84.3 212.1 ;
        RECT  78.9 206.4 81.0 207.3 ;
        RECT  84.3 206.4 88.5 207.3 ;
        RECT  80.7 202.65 81.9 203.85 ;
        RECT  83.1 202.65 84.3 203.85 ;
        RECT  80.7 211.95 81.9 213.15 ;
        RECT  83.1 211.95 84.3 213.15 ;
        RECT  85.5 211.95 86.7 213.15 ;
        RECT  85.5 201.45 86.7 202.65 ;
        RECT  81.0 206.25 82.2 207.45 ;
        RECT  66.9 208.8 68.1 210.0 ;
        RECT  51.0 208.8 52.2 210.0 ;
        RECT  50.7 229.05 51.9 230.25 ;
        RECT  57.0 229.05 58.2 230.25 ;
        RECT  57.3 229.05 66.9 229.95 ;
        RECT  57.3 214.35 66.9 215.25 ;
        RECT  63.9 215.25 65.1 217.65 ;
        RECT  63.9 227.25 65.1 229.05 ;
        RECT  59.1 228.15 60.3 229.05 ;
        RECT  59.1 215.25 60.3 216.45 ;
        RECT  61.5 217.5 62.7 226.95 ;
        RECT  57.3 222.3 59.4 223.2 ;
        RECT  62.7 222.3 66.9 223.2 ;
        RECT  59.1 223.35 60.3 224.55 ;
        RECT  61.5 223.35 62.7 224.55 ;
        RECT  59.1 222.45 60.3 223.65 ;
        RECT  61.5 222.45 62.7 223.65 ;
        RECT  63.9 217.65 65.1 218.85 ;
        RECT  63.9 228.15 65.1 229.35 ;
        RECT  59.4 223.35 60.6 224.55 ;
        RECT  66.9 229.05 78.9 229.95 ;
        RECT  66.9 214.35 78.9 215.25 ;
        RECT  75.9 214.8 76.8 217.65 ;
        RECT  75.9 227.1 76.8 229.5 ;
        RECT  68.85 214.8 69.75 217.65 ;
        RECT  73.65 214.8 74.55 217.65 ;
        RECT  68.85 226.65 69.75 229.5 ;
        RECT  66.9 219.9 69.0 220.8 ;
        RECT  66.9 223.2 72.0 224.1 ;
        RECT  74.55 222.3 78.9 223.2 ;
        RECT  68.7 221.85 69.9 223.05 ;
        RECT  71.1 221.85 72.3 223.05 ;
        RECT  71.1 221.85 72.3 223.05 ;
        RECT  73.5 221.85 74.7 223.05 ;
        RECT  68.7 222.45 69.9 223.65 ;
        RECT  71.1 222.45 72.3 223.65 ;
        RECT  71.1 222.45 72.3 223.65 ;
        RECT  73.5 222.45 74.7 223.65 ;
        RECT  75.9 217.65 77.1 218.85 ;
        RECT  75.9 227.85 77.1 229.05 ;
        RECT  74.1 234.9 75.0 235.8 ;
        RECT  71.1 234.9 72.0 235.8 ;
        RECT  74.1 227.85 75.0 235.35 ;
        RECT  71.55 234.9 74.55 235.8 ;
        RECT  71.1 235.35 72.0 238.05 ;
        RECT  69.0 221.1 70.2 222.3 ;
        RECT  72.0 224.4 73.2 225.6 ;
        RECT  78.9 229.05 88.5 229.95 ;
        RECT  78.9 214.35 88.5 215.25 ;
        RECT  85.5 215.25 86.7 217.65 ;
        RECT  85.5 227.25 86.7 229.05 ;
        RECT  80.7 228.15 81.9 229.05 ;
        RECT  80.7 215.25 81.9 216.45 ;
        RECT  83.1 217.5 84.3 226.95 ;
        RECT  78.9 222.3 81.0 223.2 ;
        RECT  84.3 222.3 88.5 223.2 ;
        RECT  80.7 223.35 81.9 224.55 ;
        RECT  83.1 223.35 84.3 224.55 ;
        RECT  80.7 222.45 81.9 223.65 ;
        RECT  83.1 222.45 84.3 223.65 ;
        RECT  85.5 217.65 86.7 218.85 ;
        RECT  85.5 228.15 86.7 229.35 ;
        RECT  81.0 223.35 82.2 224.55 ;
        RECT  66.9 219.6 68.1 220.8 ;
        RECT  51.0 219.6 52.2 220.8 ;
        RECT  50.7 243.75 51.9 244.95 ;
        RECT  57.0 243.75 58.2 244.95 ;
        RECT  57.3 229.05 66.9 229.95 ;
        RECT  57.3 243.75 66.9 244.65 ;
        RECT  63.9 241.35 65.1 243.75 ;
        RECT  63.9 229.95 65.1 231.75 ;
        RECT  59.1 229.95 60.3 230.85 ;
        RECT  59.1 242.55 60.3 243.75 ;
        RECT  61.5 232.05 62.7 241.5 ;
        RECT  57.3 235.8 59.4 236.7 ;
        RECT  62.7 235.8 66.9 236.7 ;
        RECT  59.1 232.05 60.3 233.25 ;
        RECT  61.5 232.05 62.7 233.25 ;
        RECT  59.1 241.35 60.3 242.55 ;
        RECT  61.5 241.35 62.7 242.55 ;
        RECT  63.9 241.35 65.1 242.55 ;
        RECT  63.9 230.85 65.1 232.05 ;
        RECT  59.4 235.65 60.6 236.85 ;
        RECT  66.9 229.05 78.9 229.95 ;
        RECT  66.9 243.75 78.9 244.65 ;
        RECT  75.9 241.35 76.8 244.2 ;
        RECT  75.9 229.5 76.8 231.9 ;
        RECT  68.85 241.35 69.75 244.2 ;
        RECT  73.65 241.35 74.55 244.2 ;
        RECT  68.85 229.5 69.75 232.35 ;
        RECT  66.9 238.2 69.0 239.1 ;
        RECT  66.9 234.9 72.0 235.8 ;
        RECT  74.55 235.8 78.9 236.7 ;
        RECT  68.7 232.35 69.9 233.55 ;
        RECT  71.1 232.35 72.3 233.55 ;
        RECT  71.1 232.35 72.3 233.55 ;
        RECT  73.5 232.35 74.7 233.55 ;
        RECT  68.7 241.35 69.9 242.55 ;
        RECT  71.1 241.35 72.3 242.55 ;
        RECT  71.1 241.35 72.3 242.55 ;
        RECT  73.5 241.35 74.7 242.55 ;
        RECT  75.9 241.35 77.1 242.55 ;
        RECT  75.9 231.15 77.1 232.35 ;
        RECT  74.1 238.2 75.0 239.1 ;
        RECT  71.1 238.2 72.0 239.1 ;
        RECT  74.1 231.15 75.0 238.65 ;
        RECT  71.55 238.2 74.55 239.1 ;
        RECT  71.1 238.65 72.0 241.35 ;
        RECT  69.0 237.9 70.2 239.1 ;
        RECT  72.0 234.6 73.2 235.8 ;
        RECT  78.9 229.05 88.5 229.95 ;
        RECT  78.9 243.75 88.5 244.65 ;
        RECT  85.5 241.35 86.7 243.75 ;
        RECT  85.5 229.95 86.7 231.75 ;
        RECT  80.7 229.95 81.9 230.85 ;
        RECT  80.7 242.55 81.9 243.75 ;
        RECT  83.1 232.05 84.3 241.5 ;
        RECT  78.9 235.8 81.0 236.7 ;
        RECT  84.3 235.8 88.5 236.7 ;
        RECT  80.7 232.05 81.9 233.25 ;
        RECT  83.1 232.05 84.3 233.25 ;
        RECT  80.7 241.35 81.9 242.55 ;
        RECT  83.1 241.35 84.3 242.55 ;
        RECT  85.5 241.35 86.7 242.55 ;
        RECT  85.5 230.85 86.7 232.05 ;
        RECT  81.0 235.65 82.2 236.85 ;
        RECT  66.9 238.2 68.1 239.4 ;
        RECT  51.0 238.2 52.2 239.4 ;
        RECT  50.7 258.45 51.9 259.65 ;
        RECT  57.0 258.45 58.2 259.65 ;
        RECT  57.3 258.45 66.9 259.35 ;
        RECT  57.3 243.75 66.9 244.65 ;
        RECT  63.9 244.65 65.1 247.05 ;
        RECT  63.9 256.65 65.1 258.45 ;
        RECT  59.1 257.55 60.3 258.45 ;
        RECT  59.1 244.65 60.3 245.85 ;
        RECT  61.5 246.9 62.7 256.35 ;
        RECT  57.3 251.7 59.4 252.6 ;
        RECT  62.7 251.7 66.9 252.6 ;
        RECT  59.1 252.75 60.3 253.95 ;
        RECT  61.5 252.75 62.7 253.95 ;
        RECT  59.1 251.85 60.3 253.05 ;
        RECT  61.5 251.85 62.7 253.05 ;
        RECT  63.9 247.05 65.1 248.25 ;
        RECT  63.9 257.55 65.1 258.75 ;
        RECT  59.4 252.75 60.6 253.95 ;
        RECT  66.9 258.45 78.9 259.35 ;
        RECT  66.9 243.75 78.9 244.65 ;
        RECT  75.9 244.2 76.8 247.05 ;
        RECT  75.9 256.5 76.8 258.9 ;
        RECT  68.85 244.2 69.75 247.05 ;
        RECT  73.65 244.2 74.55 247.05 ;
        RECT  68.85 256.05 69.75 258.9 ;
        RECT  66.9 249.3 69.0 250.2 ;
        RECT  66.9 252.6 72.0 253.5 ;
        RECT  74.55 251.7 78.9 252.6 ;
        RECT  68.7 251.25 69.9 252.45 ;
        RECT  71.1 251.25 72.3 252.45 ;
        RECT  71.1 251.25 72.3 252.45 ;
        RECT  73.5 251.25 74.7 252.45 ;
        RECT  68.7 251.85 69.9 253.05 ;
        RECT  71.1 251.85 72.3 253.05 ;
        RECT  71.1 251.85 72.3 253.05 ;
        RECT  73.5 251.85 74.7 253.05 ;
        RECT  75.9 247.05 77.1 248.25 ;
        RECT  75.9 257.25 77.1 258.45 ;
        RECT  74.1 264.3 75.0 265.2 ;
        RECT  71.1 264.3 72.0 265.2 ;
        RECT  74.1 257.25 75.0 264.75 ;
        RECT  71.55 264.3 74.55 265.2 ;
        RECT  71.1 264.75 72.0 267.45 ;
        RECT  69.0 250.5 70.2 251.7 ;
        RECT  72.0 253.8 73.2 255.0 ;
        RECT  78.9 258.45 88.5 259.35 ;
        RECT  78.9 243.75 88.5 244.65 ;
        RECT  85.5 244.65 86.7 247.05 ;
        RECT  85.5 256.65 86.7 258.45 ;
        RECT  80.7 257.55 81.9 258.45 ;
        RECT  80.7 244.65 81.9 245.85 ;
        RECT  83.1 246.9 84.3 256.35 ;
        RECT  78.9 251.7 81.0 252.6 ;
        RECT  84.3 251.7 88.5 252.6 ;
        RECT  80.7 252.75 81.9 253.95 ;
        RECT  83.1 252.75 84.3 253.95 ;
        RECT  80.7 251.85 81.9 253.05 ;
        RECT  83.1 251.85 84.3 253.05 ;
        RECT  85.5 247.05 86.7 248.25 ;
        RECT  85.5 257.55 86.7 258.75 ;
        RECT  81.0 252.75 82.2 253.95 ;
        RECT  66.9 249.0 68.1 250.2 ;
        RECT  51.0 249.0 52.2 250.2 ;
        RECT  50.7 273.15 51.9 274.35 ;
        RECT  57.0 273.15 58.2 274.35 ;
        RECT  57.3 258.45 66.9 259.35 ;
        RECT  57.3 273.15 66.9 274.05 ;
        RECT  63.9 270.75 65.1 273.15 ;
        RECT  63.9 259.35 65.1 261.15 ;
        RECT  59.1 259.35 60.3 260.25 ;
        RECT  59.1 271.95 60.3 273.15 ;
        RECT  61.5 261.45 62.7 270.9 ;
        RECT  57.3 265.2 59.4 266.1 ;
        RECT  62.7 265.2 66.9 266.1 ;
        RECT  59.1 261.45 60.3 262.65 ;
        RECT  61.5 261.45 62.7 262.65 ;
        RECT  59.1 270.75 60.3 271.95 ;
        RECT  61.5 270.75 62.7 271.95 ;
        RECT  63.9 270.75 65.1 271.95 ;
        RECT  63.9 260.25 65.1 261.45 ;
        RECT  59.4 265.05 60.6 266.25 ;
        RECT  66.9 258.45 78.9 259.35 ;
        RECT  66.9 273.15 78.9 274.05 ;
        RECT  75.9 270.75 76.8 273.6 ;
        RECT  75.9 258.9 76.8 261.3 ;
        RECT  68.85 270.75 69.75 273.6 ;
        RECT  73.65 270.75 74.55 273.6 ;
        RECT  68.85 258.9 69.75 261.75 ;
        RECT  66.9 267.6 69.0 268.5 ;
        RECT  66.9 264.3 72.0 265.2 ;
        RECT  74.55 265.2 78.9 266.1 ;
        RECT  68.7 261.75 69.9 262.95 ;
        RECT  71.1 261.75 72.3 262.95 ;
        RECT  71.1 261.75 72.3 262.95 ;
        RECT  73.5 261.75 74.7 262.95 ;
        RECT  68.7 270.75 69.9 271.95 ;
        RECT  71.1 270.75 72.3 271.95 ;
        RECT  71.1 270.75 72.3 271.95 ;
        RECT  73.5 270.75 74.7 271.95 ;
        RECT  75.9 270.75 77.1 271.95 ;
        RECT  75.9 260.55 77.1 261.75 ;
        RECT  74.1 267.6 75.0 268.5 ;
        RECT  71.1 267.6 72.0 268.5 ;
        RECT  74.1 260.55 75.0 268.05 ;
        RECT  71.55 267.6 74.55 268.5 ;
        RECT  71.1 268.05 72.0 270.75 ;
        RECT  69.0 267.3 70.2 268.5 ;
        RECT  72.0 264.0 73.2 265.2 ;
        RECT  78.9 258.45 88.5 259.35 ;
        RECT  78.9 273.15 88.5 274.05 ;
        RECT  85.5 270.75 86.7 273.15 ;
        RECT  85.5 259.35 86.7 261.15 ;
        RECT  80.7 259.35 81.9 260.25 ;
        RECT  80.7 271.95 81.9 273.15 ;
        RECT  83.1 261.45 84.3 270.9 ;
        RECT  78.9 265.2 81.0 266.1 ;
        RECT  84.3 265.2 88.5 266.1 ;
        RECT  80.7 261.45 81.9 262.65 ;
        RECT  83.1 261.45 84.3 262.65 ;
        RECT  80.7 270.75 81.9 271.95 ;
        RECT  83.1 270.75 84.3 271.95 ;
        RECT  85.5 270.75 86.7 271.95 ;
        RECT  85.5 260.25 86.7 261.45 ;
        RECT  81.0 265.05 82.2 266.25 ;
        RECT  66.9 267.6 68.1 268.8 ;
        RECT  51.0 267.6 52.2 268.8 ;
        RECT  50.7 287.85 51.9 289.05 ;
        RECT  57.0 287.85 58.2 289.05 ;
        RECT  57.3 287.85 66.9 288.75 ;
        RECT  57.3 273.15 66.9 274.05 ;
        RECT  63.9 274.05 65.1 276.45 ;
        RECT  63.9 286.05 65.1 287.85 ;
        RECT  59.1 286.95 60.3 287.85 ;
        RECT  59.1 274.05 60.3 275.25 ;
        RECT  61.5 276.3 62.7 285.75 ;
        RECT  57.3 281.1 59.4 282.0 ;
        RECT  62.7 281.1 66.9 282.0 ;
        RECT  59.1 282.15 60.3 283.35 ;
        RECT  61.5 282.15 62.7 283.35 ;
        RECT  59.1 281.25 60.3 282.45 ;
        RECT  61.5 281.25 62.7 282.45 ;
        RECT  63.9 276.45 65.1 277.65 ;
        RECT  63.9 286.95 65.1 288.15 ;
        RECT  59.4 282.15 60.6 283.35 ;
        RECT  66.9 287.85 78.9 288.75 ;
        RECT  66.9 273.15 78.9 274.05 ;
        RECT  75.9 273.6 76.8 276.45 ;
        RECT  75.9 285.9 76.8 288.3 ;
        RECT  68.85 273.6 69.75 276.45 ;
        RECT  73.65 273.6 74.55 276.45 ;
        RECT  68.85 285.45 69.75 288.3 ;
        RECT  66.9 278.7 69.0 279.6 ;
        RECT  66.9 282.0 72.0 282.9 ;
        RECT  74.55 281.1 78.9 282.0 ;
        RECT  68.7 280.65 69.9 281.85 ;
        RECT  71.1 280.65 72.3 281.85 ;
        RECT  71.1 280.65 72.3 281.85 ;
        RECT  73.5 280.65 74.7 281.85 ;
        RECT  68.7 281.25 69.9 282.45 ;
        RECT  71.1 281.25 72.3 282.45 ;
        RECT  71.1 281.25 72.3 282.45 ;
        RECT  73.5 281.25 74.7 282.45 ;
        RECT  75.9 276.45 77.1 277.65 ;
        RECT  75.9 286.65 77.1 287.85 ;
        RECT  74.1 293.7 75.0 294.6 ;
        RECT  71.1 293.7 72.0 294.6 ;
        RECT  74.1 286.65 75.0 294.15 ;
        RECT  71.55 293.7 74.55 294.6 ;
        RECT  71.1 294.15 72.0 296.85 ;
        RECT  69.0 279.9 70.2 281.1 ;
        RECT  72.0 283.2 73.2 284.4 ;
        RECT  78.9 287.85 88.5 288.75 ;
        RECT  78.9 273.15 88.5 274.05 ;
        RECT  85.5 274.05 86.7 276.45 ;
        RECT  85.5 286.05 86.7 287.85 ;
        RECT  80.7 286.95 81.9 287.85 ;
        RECT  80.7 274.05 81.9 275.25 ;
        RECT  83.1 276.3 84.3 285.75 ;
        RECT  78.9 281.1 81.0 282.0 ;
        RECT  84.3 281.1 88.5 282.0 ;
        RECT  80.7 282.15 81.9 283.35 ;
        RECT  83.1 282.15 84.3 283.35 ;
        RECT  80.7 281.25 81.9 282.45 ;
        RECT  83.1 281.25 84.3 282.45 ;
        RECT  85.5 276.45 86.7 277.65 ;
        RECT  85.5 286.95 86.7 288.15 ;
        RECT  81.0 282.15 82.2 283.35 ;
        RECT  66.9 278.4 68.1 279.6 ;
        RECT  51.0 278.4 52.2 279.6 ;
        RECT  50.7 302.55 51.9 303.75 ;
        RECT  57.0 302.55 58.2 303.75 ;
        RECT  57.3 287.85 66.9 288.75 ;
        RECT  57.3 302.55 66.9 303.45 ;
        RECT  63.9 300.15 65.1 302.55 ;
        RECT  63.9 288.75 65.1 290.55 ;
        RECT  59.1 288.75 60.3 289.65 ;
        RECT  59.1 301.35 60.3 302.55 ;
        RECT  61.5 290.85 62.7 300.3 ;
        RECT  57.3 294.6 59.4 295.5 ;
        RECT  62.7 294.6 66.9 295.5 ;
        RECT  59.1 290.85 60.3 292.05 ;
        RECT  61.5 290.85 62.7 292.05 ;
        RECT  59.1 300.15 60.3 301.35 ;
        RECT  61.5 300.15 62.7 301.35 ;
        RECT  63.9 300.15 65.1 301.35 ;
        RECT  63.9 289.65 65.1 290.85 ;
        RECT  59.4 294.45 60.6 295.65 ;
        RECT  66.9 287.85 78.9 288.75 ;
        RECT  66.9 302.55 78.9 303.45 ;
        RECT  75.9 300.15 76.8 303.0 ;
        RECT  75.9 288.3 76.8 290.7 ;
        RECT  68.85 300.15 69.75 303.0 ;
        RECT  73.65 300.15 74.55 303.0 ;
        RECT  68.85 288.3 69.75 291.15 ;
        RECT  66.9 297.0 69.0 297.9 ;
        RECT  66.9 293.7 72.0 294.6 ;
        RECT  74.55 294.6 78.9 295.5 ;
        RECT  68.7 291.15 69.9 292.35 ;
        RECT  71.1 291.15 72.3 292.35 ;
        RECT  71.1 291.15 72.3 292.35 ;
        RECT  73.5 291.15 74.7 292.35 ;
        RECT  68.7 300.15 69.9 301.35 ;
        RECT  71.1 300.15 72.3 301.35 ;
        RECT  71.1 300.15 72.3 301.35 ;
        RECT  73.5 300.15 74.7 301.35 ;
        RECT  75.9 300.15 77.1 301.35 ;
        RECT  75.9 289.95 77.1 291.15 ;
        RECT  74.1 297.0 75.0 297.9 ;
        RECT  71.1 297.0 72.0 297.9 ;
        RECT  74.1 289.95 75.0 297.45 ;
        RECT  71.55 297.0 74.55 297.9 ;
        RECT  71.1 297.45 72.0 300.15 ;
        RECT  69.0 296.7 70.2 297.9 ;
        RECT  72.0 293.4 73.2 294.6 ;
        RECT  78.9 287.85 88.5 288.75 ;
        RECT  78.9 302.55 88.5 303.45 ;
        RECT  85.5 300.15 86.7 302.55 ;
        RECT  85.5 288.75 86.7 290.55 ;
        RECT  80.7 288.75 81.9 289.65 ;
        RECT  80.7 301.35 81.9 302.55 ;
        RECT  83.1 290.85 84.3 300.3 ;
        RECT  78.9 294.6 81.0 295.5 ;
        RECT  84.3 294.6 88.5 295.5 ;
        RECT  80.7 290.85 81.9 292.05 ;
        RECT  83.1 290.85 84.3 292.05 ;
        RECT  80.7 300.15 81.9 301.35 ;
        RECT  83.1 300.15 84.3 301.35 ;
        RECT  85.5 300.15 86.7 301.35 ;
        RECT  85.5 289.65 86.7 290.85 ;
        RECT  81.0 294.45 82.2 295.65 ;
        RECT  66.9 297.0 68.1 298.2 ;
        RECT  51.0 297.0 52.2 298.2 ;
        RECT  50.7 317.25 51.9 318.45 ;
        RECT  57.0 317.25 58.2 318.45 ;
        RECT  57.3 317.25 66.9 318.15 ;
        RECT  57.3 302.55 66.9 303.45 ;
        RECT  63.9 303.45 65.1 305.85 ;
        RECT  63.9 315.45 65.1 317.25 ;
        RECT  59.1 316.35 60.3 317.25 ;
        RECT  59.1 303.45 60.3 304.65 ;
        RECT  61.5 305.7 62.7 315.15 ;
        RECT  57.3 310.5 59.4 311.4 ;
        RECT  62.7 310.5 66.9 311.4 ;
        RECT  59.1 311.55 60.3 312.75 ;
        RECT  61.5 311.55 62.7 312.75 ;
        RECT  59.1 310.65 60.3 311.85 ;
        RECT  61.5 310.65 62.7 311.85 ;
        RECT  63.9 305.85 65.1 307.05 ;
        RECT  63.9 316.35 65.1 317.55 ;
        RECT  59.4 311.55 60.6 312.75 ;
        RECT  66.9 317.25 78.9 318.15 ;
        RECT  66.9 302.55 78.9 303.45 ;
        RECT  75.9 303.0 76.8 305.85 ;
        RECT  75.9 315.3 76.8 317.7 ;
        RECT  68.85 303.0 69.75 305.85 ;
        RECT  73.65 303.0 74.55 305.85 ;
        RECT  68.85 314.85 69.75 317.7 ;
        RECT  66.9 308.1 69.0 309.0 ;
        RECT  66.9 311.4 72.0 312.3 ;
        RECT  74.55 310.5 78.9 311.4 ;
        RECT  68.7 310.05 69.9 311.25 ;
        RECT  71.1 310.05 72.3 311.25 ;
        RECT  71.1 310.05 72.3 311.25 ;
        RECT  73.5 310.05 74.7 311.25 ;
        RECT  68.7 310.65 69.9 311.85 ;
        RECT  71.1 310.65 72.3 311.85 ;
        RECT  71.1 310.65 72.3 311.85 ;
        RECT  73.5 310.65 74.7 311.85 ;
        RECT  75.9 305.85 77.1 307.05 ;
        RECT  75.9 316.05 77.1 317.25 ;
        RECT  74.1 323.1 75.0 324.0 ;
        RECT  71.1 323.1 72.0 324.0 ;
        RECT  74.1 316.05 75.0 323.55 ;
        RECT  71.55 323.1 74.55 324.0 ;
        RECT  71.1 323.55 72.0 326.25 ;
        RECT  69.0 309.3 70.2 310.5 ;
        RECT  72.0 312.6 73.2 313.8 ;
        RECT  78.9 317.25 88.5 318.15 ;
        RECT  78.9 302.55 88.5 303.45 ;
        RECT  85.5 303.45 86.7 305.85 ;
        RECT  85.5 315.45 86.7 317.25 ;
        RECT  80.7 316.35 81.9 317.25 ;
        RECT  80.7 303.45 81.9 304.65 ;
        RECT  83.1 305.7 84.3 315.15 ;
        RECT  78.9 310.5 81.0 311.4 ;
        RECT  84.3 310.5 88.5 311.4 ;
        RECT  80.7 311.55 81.9 312.75 ;
        RECT  83.1 311.55 84.3 312.75 ;
        RECT  80.7 310.65 81.9 311.85 ;
        RECT  83.1 310.65 84.3 311.85 ;
        RECT  85.5 305.85 86.7 307.05 ;
        RECT  85.5 316.35 86.7 317.55 ;
        RECT  81.0 311.55 82.2 312.75 ;
        RECT  66.9 307.8 68.1 309.0 ;
        RECT  51.0 307.8 52.2 309.0 ;
        RECT  50.7 331.95 51.9 333.15 ;
        RECT  57.0 331.95 58.2 333.15 ;
        RECT  57.3 317.25 66.9 318.15 ;
        RECT  57.3 331.95 66.9 332.85 ;
        RECT  63.9 329.55 65.1 331.95 ;
        RECT  63.9 318.15 65.1 319.95 ;
        RECT  59.1 318.15 60.3 319.05 ;
        RECT  59.1 330.75 60.3 331.95 ;
        RECT  61.5 320.25 62.7 329.7 ;
        RECT  57.3 324.0 59.4 324.9 ;
        RECT  62.7 324.0 66.9 324.9 ;
        RECT  59.1 320.25 60.3 321.45 ;
        RECT  61.5 320.25 62.7 321.45 ;
        RECT  59.1 329.55 60.3 330.75 ;
        RECT  61.5 329.55 62.7 330.75 ;
        RECT  63.9 329.55 65.1 330.75 ;
        RECT  63.9 319.05 65.1 320.25 ;
        RECT  59.4 323.85 60.6 325.05 ;
        RECT  66.9 317.25 78.9 318.15 ;
        RECT  66.9 331.95 78.9 332.85 ;
        RECT  75.9 329.55 76.8 332.4 ;
        RECT  75.9 317.7 76.8 320.1 ;
        RECT  68.85 329.55 69.75 332.4 ;
        RECT  73.65 329.55 74.55 332.4 ;
        RECT  68.85 317.7 69.75 320.55 ;
        RECT  66.9 326.4 69.0 327.3 ;
        RECT  66.9 323.1 72.0 324.0 ;
        RECT  74.55 324.0 78.9 324.9 ;
        RECT  68.7 320.55 69.9 321.75 ;
        RECT  71.1 320.55 72.3 321.75 ;
        RECT  71.1 320.55 72.3 321.75 ;
        RECT  73.5 320.55 74.7 321.75 ;
        RECT  68.7 329.55 69.9 330.75 ;
        RECT  71.1 329.55 72.3 330.75 ;
        RECT  71.1 329.55 72.3 330.75 ;
        RECT  73.5 329.55 74.7 330.75 ;
        RECT  75.9 329.55 77.1 330.75 ;
        RECT  75.9 319.35 77.1 320.55 ;
        RECT  74.1 326.4 75.0 327.3 ;
        RECT  71.1 326.4 72.0 327.3 ;
        RECT  74.1 319.35 75.0 326.85 ;
        RECT  71.55 326.4 74.55 327.3 ;
        RECT  71.1 326.85 72.0 329.55 ;
        RECT  69.0 326.1 70.2 327.3 ;
        RECT  72.0 322.8 73.2 324.0 ;
        RECT  78.9 317.25 88.5 318.15 ;
        RECT  78.9 331.95 88.5 332.85 ;
        RECT  85.5 329.55 86.7 331.95 ;
        RECT  85.5 318.15 86.7 319.95 ;
        RECT  80.7 318.15 81.9 319.05 ;
        RECT  80.7 330.75 81.9 331.95 ;
        RECT  83.1 320.25 84.3 329.7 ;
        RECT  78.9 324.0 81.0 324.9 ;
        RECT  84.3 324.0 88.5 324.9 ;
        RECT  80.7 320.25 81.9 321.45 ;
        RECT  83.1 320.25 84.3 321.45 ;
        RECT  80.7 329.55 81.9 330.75 ;
        RECT  83.1 329.55 84.3 330.75 ;
        RECT  85.5 329.55 86.7 330.75 ;
        RECT  85.5 319.05 86.7 320.25 ;
        RECT  81.0 323.85 82.2 325.05 ;
        RECT  66.9 326.4 68.1 327.6 ;
        RECT  51.0 326.4 52.2 327.6 ;
        RECT  50.7 346.65 51.9 347.85 ;
        RECT  57.0 346.65 58.2 347.85 ;
        RECT  57.3 346.65 66.9 347.55 ;
        RECT  57.3 331.95 66.9 332.85 ;
        RECT  63.9 332.85 65.1 335.25 ;
        RECT  63.9 344.85 65.1 346.65 ;
        RECT  59.1 345.75 60.3 346.65 ;
        RECT  59.1 332.85 60.3 334.05 ;
        RECT  61.5 335.1 62.7 344.55 ;
        RECT  57.3 339.9 59.4 340.8 ;
        RECT  62.7 339.9 66.9 340.8 ;
        RECT  59.1 340.95 60.3 342.15 ;
        RECT  61.5 340.95 62.7 342.15 ;
        RECT  59.1 340.05 60.3 341.25 ;
        RECT  61.5 340.05 62.7 341.25 ;
        RECT  63.9 335.25 65.1 336.45 ;
        RECT  63.9 345.75 65.1 346.95 ;
        RECT  59.4 340.95 60.6 342.15 ;
        RECT  66.9 346.65 78.9 347.55 ;
        RECT  66.9 331.95 78.9 332.85 ;
        RECT  75.9 332.4 76.8 335.25 ;
        RECT  75.9 344.7 76.8 347.1 ;
        RECT  68.85 332.4 69.75 335.25 ;
        RECT  73.65 332.4 74.55 335.25 ;
        RECT  68.85 344.25 69.75 347.1 ;
        RECT  66.9 337.5 69.0 338.4 ;
        RECT  66.9 340.8 72.0 341.7 ;
        RECT  74.55 339.9 78.9 340.8 ;
        RECT  68.7 339.45 69.9 340.65 ;
        RECT  71.1 339.45 72.3 340.65 ;
        RECT  71.1 339.45 72.3 340.65 ;
        RECT  73.5 339.45 74.7 340.65 ;
        RECT  68.7 340.05 69.9 341.25 ;
        RECT  71.1 340.05 72.3 341.25 ;
        RECT  71.1 340.05 72.3 341.25 ;
        RECT  73.5 340.05 74.7 341.25 ;
        RECT  75.9 335.25 77.1 336.45 ;
        RECT  75.9 345.45 77.1 346.65 ;
        RECT  74.1 352.5 75.0 353.4 ;
        RECT  71.1 352.5 72.0 353.4 ;
        RECT  74.1 345.45 75.0 352.95 ;
        RECT  71.55 352.5 74.55 353.4 ;
        RECT  71.1 352.95 72.0 355.65 ;
        RECT  69.0 338.7 70.2 339.9 ;
        RECT  72.0 342.0 73.2 343.2 ;
        RECT  78.9 346.65 88.5 347.55 ;
        RECT  78.9 331.95 88.5 332.85 ;
        RECT  85.5 332.85 86.7 335.25 ;
        RECT  85.5 344.85 86.7 346.65 ;
        RECT  80.7 345.75 81.9 346.65 ;
        RECT  80.7 332.85 81.9 334.05 ;
        RECT  83.1 335.1 84.3 344.55 ;
        RECT  78.9 339.9 81.0 340.8 ;
        RECT  84.3 339.9 88.5 340.8 ;
        RECT  80.7 340.95 81.9 342.15 ;
        RECT  83.1 340.95 84.3 342.15 ;
        RECT  80.7 340.05 81.9 341.25 ;
        RECT  83.1 340.05 84.3 341.25 ;
        RECT  85.5 335.25 86.7 336.45 ;
        RECT  85.5 345.75 86.7 346.95 ;
        RECT  81.0 340.95 82.2 342.15 ;
        RECT  66.9 337.2 68.1 338.4 ;
        RECT  51.0 337.2 52.2 338.4 ;
        RECT  50.7 361.35 51.9 362.55 ;
        RECT  57.0 361.35 58.2 362.55 ;
        RECT  57.3 346.65 66.9 347.55 ;
        RECT  57.3 361.35 66.9 362.25 ;
        RECT  63.9 358.95 65.1 361.35 ;
        RECT  63.9 347.55 65.1 349.35 ;
        RECT  59.1 347.55 60.3 348.45 ;
        RECT  59.1 360.15 60.3 361.35 ;
        RECT  61.5 349.65 62.7 359.1 ;
        RECT  57.3 353.4 59.4 354.3 ;
        RECT  62.7 353.4 66.9 354.3 ;
        RECT  59.1 349.65 60.3 350.85 ;
        RECT  61.5 349.65 62.7 350.85 ;
        RECT  59.1 358.95 60.3 360.15 ;
        RECT  61.5 358.95 62.7 360.15 ;
        RECT  63.9 358.95 65.1 360.15 ;
        RECT  63.9 348.45 65.1 349.65 ;
        RECT  59.4 353.25 60.6 354.45 ;
        RECT  66.9 346.65 78.9 347.55 ;
        RECT  66.9 361.35 78.9 362.25 ;
        RECT  75.9 358.95 76.8 361.8 ;
        RECT  75.9 347.1 76.8 349.5 ;
        RECT  68.85 358.95 69.75 361.8 ;
        RECT  73.65 358.95 74.55 361.8 ;
        RECT  68.85 347.1 69.75 349.95 ;
        RECT  66.9 355.8 69.0 356.7 ;
        RECT  66.9 352.5 72.0 353.4 ;
        RECT  74.55 353.4 78.9 354.3 ;
        RECT  68.7 349.95 69.9 351.15 ;
        RECT  71.1 349.95 72.3 351.15 ;
        RECT  71.1 349.95 72.3 351.15 ;
        RECT  73.5 349.95 74.7 351.15 ;
        RECT  68.7 358.95 69.9 360.15 ;
        RECT  71.1 358.95 72.3 360.15 ;
        RECT  71.1 358.95 72.3 360.15 ;
        RECT  73.5 358.95 74.7 360.15 ;
        RECT  75.9 358.95 77.1 360.15 ;
        RECT  75.9 348.75 77.1 349.95 ;
        RECT  74.1 355.8 75.0 356.7 ;
        RECT  71.1 355.8 72.0 356.7 ;
        RECT  74.1 348.75 75.0 356.25 ;
        RECT  71.55 355.8 74.55 356.7 ;
        RECT  71.1 356.25 72.0 358.95 ;
        RECT  69.0 355.5 70.2 356.7 ;
        RECT  72.0 352.2 73.2 353.4 ;
        RECT  78.9 346.65 88.5 347.55 ;
        RECT  78.9 361.35 88.5 362.25 ;
        RECT  85.5 358.95 86.7 361.35 ;
        RECT  85.5 347.55 86.7 349.35 ;
        RECT  80.7 347.55 81.9 348.45 ;
        RECT  80.7 360.15 81.9 361.35 ;
        RECT  83.1 349.65 84.3 359.1 ;
        RECT  78.9 353.4 81.0 354.3 ;
        RECT  84.3 353.4 88.5 354.3 ;
        RECT  80.7 349.65 81.9 350.85 ;
        RECT  83.1 349.65 84.3 350.85 ;
        RECT  80.7 358.95 81.9 360.15 ;
        RECT  83.1 358.95 84.3 360.15 ;
        RECT  85.5 358.95 86.7 360.15 ;
        RECT  85.5 348.45 86.7 349.65 ;
        RECT  81.0 353.25 82.2 354.45 ;
        RECT  66.9 355.8 68.1 357.0 ;
        RECT  51.0 355.8 52.2 357.0 ;
        RECT  50.7 376.05 51.9 377.25 ;
        RECT  57.0 376.05 58.2 377.25 ;
        RECT  57.3 376.05 66.9 376.95 ;
        RECT  57.3 361.35 66.9 362.25 ;
        RECT  63.9 362.25 65.1 364.65 ;
        RECT  63.9 374.25 65.1 376.05 ;
        RECT  59.1 375.15 60.3 376.05 ;
        RECT  59.1 362.25 60.3 363.45 ;
        RECT  61.5 364.5 62.7 373.95 ;
        RECT  57.3 369.3 59.4 370.2 ;
        RECT  62.7 369.3 66.9 370.2 ;
        RECT  59.1 370.35 60.3 371.55 ;
        RECT  61.5 370.35 62.7 371.55 ;
        RECT  59.1 369.45 60.3 370.65 ;
        RECT  61.5 369.45 62.7 370.65 ;
        RECT  63.9 364.65 65.1 365.85 ;
        RECT  63.9 375.15 65.1 376.35 ;
        RECT  59.4 370.35 60.6 371.55 ;
        RECT  66.9 376.05 78.9 376.95 ;
        RECT  66.9 361.35 78.9 362.25 ;
        RECT  75.9 361.8 76.8 364.65 ;
        RECT  75.9 374.1 76.8 376.5 ;
        RECT  68.85 361.8 69.75 364.65 ;
        RECT  73.65 361.8 74.55 364.65 ;
        RECT  68.85 373.65 69.75 376.5 ;
        RECT  66.9 366.9 69.0 367.8 ;
        RECT  66.9 370.2 72.0 371.1 ;
        RECT  74.55 369.3 78.9 370.2 ;
        RECT  68.7 368.85 69.9 370.05 ;
        RECT  71.1 368.85 72.3 370.05 ;
        RECT  71.1 368.85 72.3 370.05 ;
        RECT  73.5 368.85 74.7 370.05 ;
        RECT  68.7 369.45 69.9 370.65 ;
        RECT  71.1 369.45 72.3 370.65 ;
        RECT  71.1 369.45 72.3 370.65 ;
        RECT  73.5 369.45 74.7 370.65 ;
        RECT  75.9 364.65 77.1 365.85 ;
        RECT  75.9 374.85 77.1 376.05 ;
        RECT  74.1 381.9 75.0 382.8 ;
        RECT  71.1 381.9 72.0 382.8 ;
        RECT  74.1 374.85 75.0 382.35 ;
        RECT  71.55 381.9 74.55 382.8 ;
        RECT  71.1 382.35 72.0 385.05 ;
        RECT  69.0 368.1 70.2 369.3 ;
        RECT  72.0 371.4 73.2 372.6 ;
        RECT  78.9 376.05 88.5 376.95 ;
        RECT  78.9 361.35 88.5 362.25 ;
        RECT  85.5 362.25 86.7 364.65 ;
        RECT  85.5 374.25 86.7 376.05 ;
        RECT  80.7 375.15 81.9 376.05 ;
        RECT  80.7 362.25 81.9 363.45 ;
        RECT  83.1 364.5 84.3 373.95 ;
        RECT  78.9 369.3 81.0 370.2 ;
        RECT  84.3 369.3 88.5 370.2 ;
        RECT  80.7 370.35 81.9 371.55 ;
        RECT  83.1 370.35 84.3 371.55 ;
        RECT  80.7 369.45 81.9 370.65 ;
        RECT  83.1 369.45 84.3 370.65 ;
        RECT  85.5 364.65 86.7 365.85 ;
        RECT  85.5 375.15 86.7 376.35 ;
        RECT  81.0 370.35 82.2 371.55 ;
        RECT  66.9 366.6 68.1 367.8 ;
        RECT  51.0 366.6 52.2 367.8 ;
        RECT  50.7 390.75 51.9 391.95 ;
        RECT  57.0 390.75 58.2 391.95 ;
        RECT  57.3 376.05 66.9 376.95 ;
        RECT  57.3 390.75 66.9 391.65 ;
        RECT  63.9 388.35 65.1 390.75 ;
        RECT  63.9 376.95 65.1 378.75 ;
        RECT  59.1 376.95 60.3 377.85 ;
        RECT  59.1 389.55 60.3 390.75 ;
        RECT  61.5 379.05 62.7 388.5 ;
        RECT  57.3 382.8 59.4 383.7 ;
        RECT  62.7 382.8 66.9 383.7 ;
        RECT  59.1 379.05 60.3 380.25 ;
        RECT  61.5 379.05 62.7 380.25 ;
        RECT  59.1 388.35 60.3 389.55 ;
        RECT  61.5 388.35 62.7 389.55 ;
        RECT  63.9 388.35 65.1 389.55 ;
        RECT  63.9 377.85 65.1 379.05 ;
        RECT  59.4 382.65 60.6 383.85 ;
        RECT  66.9 376.05 78.9 376.95 ;
        RECT  66.9 390.75 78.9 391.65 ;
        RECT  75.9 388.35 76.8 391.2 ;
        RECT  75.9 376.5 76.8 378.9 ;
        RECT  68.85 388.35 69.75 391.2 ;
        RECT  73.65 388.35 74.55 391.2 ;
        RECT  68.85 376.5 69.75 379.35 ;
        RECT  66.9 385.2 69.0 386.1 ;
        RECT  66.9 381.9 72.0 382.8 ;
        RECT  74.55 382.8 78.9 383.7 ;
        RECT  68.7 379.35 69.9 380.55 ;
        RECT  71.1 379.35 72.3 380.55 ;
        RECT  71.1 379.35 72.3 380.55 ;
        RECT  73.5 379.35 74.7 380.55 ;
        RECT  68.7 388.35 69.9 389.55 ;
        RECT  71.1 388.35 72.3 389.55 ;
        RECT  71.1 388.35 72.3 389.55 ;
        RECT  73.5 388.35 74.7 389.55 ;
        RECT  75.9 388.35 77.1 389.55 ;
        RECT  75.9 378.15 77.1 379.35 ;
        RECT  74.1 385.2 75.0 386.1 ;
        RECT  71.1 385.2 72.0 386.1 ;
        RECT  74.1 378.15 75.0 385.65 ;
        RECT  71.55 385.2 74.55 386.1 ;
        RECT  71.1 385.65 72.0 388.35 ;
        RECT  69.0 384.9 70.2 386.1 ;
        RECT  72.0 381.6 73.2 382.8 ;
        RECT  78.9 376.05 88.5 376.95 ;
        RECT  78.9 390.75 88.5 391.65 ;
        RECT  85.5 388.35 86.7 390.75 ;
        RECT  85.5 376.95 86.7 378.75 ;
        RECT  80.7 376.95 81.9 377.85 ;
        RECT  80.7 389.55 81.9 390.75 ;
        RECT  83.1 379.05 84.3 388.5 ;
        RECT  78.9 382.8 81.0 383.7 ;
        RECT  84.3 382.8 88.5 383.7 ;
        RECT  80.7 379.05 81.9 380.25 ;
        RECT  83.1 379.05 84.3 380.25 ;
        RECT  80.7 388.35 81.9 389.55 ;
        RECT  83.1 388.35 84.3 389.55 ;
        RECT  85.5 388.35 86.7 389.55 ;
        RECT  85.5 377.85 86.7 379.05 ;
        RECT  81.0 382.65 82.2 383.85 ;
        RECT  66.9 385.2 68.1 386.4 ;
        RECT  51.0 385.2 52.2 386.4 ;
        RECT  50.7 405.45 51.9 406.65 ;
        RECT  57.0 405.45 58.2 406.65 ;
        RECT  57.3 405.45 66.9 406.35 ;
        RECT  57.3 390.75 66.9 391.65 ;
        RECT  63.9 391.65 65.1 394.05 ;
        RECT  63.9 403.65 65.1 405.45 ;
        RECT  59.1 404.55 60.3 405.45 ;
        RECT  59.1 391.65 60.3 392.85 ;
        RECT  61.5 393.9 62.7 403.35 ;
        RECT  57.3 398.7 59.4 399.6 ;
        RECT  62.7 398.7 66.9 399.6 ;
        RECT  59.1 399.75 60.3 400.95 ;
        RECT  61.5 399.75 62.7 400.95 ;
        RECT  59.1 398.85 60.3 400.05 ;
        RECT  61.5 398.85 62.7 400.05 ;
        RECT  63.9 394.05 65.1 395.25 ;
        RECT  63.9 404.55 65.1 405.75 ;
        RECT  59.4 399.75 60.6 400.95 ;
        RECT  66.9 405.45 78.9 406.35 ;
        RECT  66.9 390.75 78.9 391.65 ;
        RECT  75.9 391.2 76.8 394.05 ;
        RECT  75.9 403.5 76.8 405.9 ;
        RECT  68.85 391.2 69.75 394.05 ;
        RECT  73.65 391.2 74.55 394.05 ;
        RECT  68.85 403.05 69.75 405.9 ;
        RECT  66.9 396.3 69.0 397.2 ;
        RECT  66.9 399.6 72.0 400.5 ;
        RECT  74.55 398.7 78.9 399.6 ;
        RECT  68.7 398.25 69.9 399.45 ;
        RECT  71.1 398.25 72.3 399.45 ;
        RECT  71.1 398.25 72.3 399.45 ;
        RECT  73.5 398.25 74.7 399.45 ;
        RECT  68.7 398.85 69.9 400.05 ;
        RECT  71.1 398.85 72.3 400.05 ;
        RECT  71.1 398.85 72.3 400.05 ;
        RECT  73.5 398.85 74.7 400.05 ;
        RECT  75.9 394.05 77.1 395.25 ;
        RECT  75.9 404.25 77.1 405.45 ;
        RECT  74.1 411.3 75.0 412.2 ;
        RECT  71.1 411.3 72.0 412.2 ;
        RECT  74.1 404.25 75.0 411.75 ;
        RECT  71.55 411.3 74.55 412.2 ;
        RECT  71.1 411.75 72.0 414.45 ;
        RECT  69.0 397.5 70.2 398.7 ;
        RECT  72.0 400.8 73.2 402.0 ;
        RECT  78.9 405.45 88.5 406.35 ;
        RECT  78.9 390.75 88.5 391.65 ;
        RECT  85.5 391.65 86.7 394.05 ;
        RECT  85.5 403.65 86.7 405.45 ;
        RECT  80.7 404.55 81.9 405.45 ;
        RECT  80.7 391.65 81.9 392.85 ;
        RECT  83.1 393.9 84.3 403.35 ;
        RECT  78.9 398.7 81.0 399.6 ;
        RECT  84.3 398.7 88.5 399.6 ;
        RECT  80.7 399.75 81.9 400.95 ;
        RECT  83.1 399.75 84.3 400.95 ;
        RECT  80.7 398.85 81.9 400.05 ;
        RECT  83.1 398.85 84.3 400.05 ;
        RECT  85.5 394.05 86.7 395.25 ;
        RECT  85.5 404.55 86.7 405.75 ;
        RECT  81.0 399.75 82.2 400.95 ;
        RECT  66.9 396.0 68.1 397.2 ;
        RECT  51.0 396.0 52.2 397.2 ;
        RECT  50.7 420.15 51.9 421.35 ;
        RECT  57.0 420.15 58.2 421.35 ;
        RECT  57.3 405.45 66.9 406.35 ;
        RECT  57.3 420.15 66.9 421.05 ;
        RECT  63.9 417.75 65.1 420.15 ;
        RECT  63.9 406.35 65.1 408.15 ;
        RECT  59.1 406.35 60.3 407.25 ;
        RECT  59.1 418.95 60.3 420.15 ;
        RECT  61.5 408.45 62.7 417.9 ;
        RECT  57.3 412.2 59.4 413.1 ;
        RECT  62.7 412.2 66.9 413.1 ;
        RECT  59.1 408.45 60.3 409.65 ;
        RECT  61.5 408.45 62.7 409.65 ;
        RECT  59.1 417.75 60.3 418.95 ;
        RECT  61.5 417.75 62.7 418.95 ;
        RECT  63.9 417.75 65.1 418.95 ;
        RECT  63.9 407.25 65.1 408.45 ;
        RECT  59.4 412.05 60.6 413.25 ;
        RECT  66.9 405.45 78.9 406.35 ;
        RECT  66.9 420.15 78.9 421.05 ;
        RECT  75.9 417.75 76.8 420.6 ;
        RECT  75.9 405.9 76.8 408.3 ;
        RECT  68.85 417.75 69.75 420.6 ;
        RECT  73.65 417.75 74.55 420.6 ;
        RECT  68.85 405.9 69.75 408.75 ;
        RECT  66.9 414.6 69.0 415.5 ;
        RECT  66.9 411.3 72.0 412.2 ;
        RECT  74.55 412.2 78.9 413.1 ;
        RECT  68.7 408.75 69.9 409.95 ;
        RECT  71.1 408.75 72.3 409.95 ;
        RECT  71.1 408.75 72.3 409.95 ;
        RECT  73.5 408.75 74.7 409.95 ;
        RECT  68.7 417.75 69.9 418.95 ;
        RECT  71.1 417.75 72.3 418.95 ;
        RECT  71.1 417.75 72.3 418.95 ;
        RECT  73.5 417.75 74.7 418.95 ;
        RECT  75.9 417.75 77.1 418.95 ;
        RECT  75.9 407.55 77.1 408.75 ;
        RECT  74.1 414.6 75.0 415.5 ;
        RECT  71.1 414.6 72.0 415.5 ;
        RECT  74.1 407.55 75.0 415.05 ;
        RECT  71.55 414.6 74.55 415.5 ;
        RECT  71.1 415.05 72.0 417.75 ;
        RECT  69.0 414.3 70.2 415.5 ;
        RECT  72.0 411.0 73.2 412.2 ;
        RECT  78.9 405.45 88.5 406.35 ;
        RECT  78.9 420.15 88.5 421.05 ;
        RECT  85.5 417.75 86.7 420.15 ;
        RECT  85.5 406.35 86.7 408.15 ;
        RECT  80.7 406.35 81.9 407.25 ;
        RECT  80.7 418.95 81.9 420.15 ;
        RECT  83.1 408.45 84.3 417.9 ;
        RECT  78.9 412.2 81.0 413.1 ;
        RECT  84.3 412.2 88.5 413.1 ;
        RECT  80.7 408.45 81.9 409.65 ;
        RECT  83.1 408.45 84.3 409.65 ;
        RECT  80.7 417.75 81.9 418.95 ;
        RECT  83.1 417.75 84.3 418.95 ;
        RECT  85.5 417.75 86.7 418.95 ;
        RECT  85.5 407.25 86.7 408.45 ;
        RECT  81.0 412.05 82.2 413.25 ;
        RECT  66.9 414.6 68.1 415.8 ;
        RECT  51.0 414.6 52.2 415.8 ;
        RECT  50.7 434.85 51.9 436.05 ;
        RECT  57.0 434.85 58.2 436.05 ;
        RECT  57.3 434.85 66.9 435.75 ;
        RECT  57.3 420.15 66.9 421.05 ;
        RECT  63.9 421.05 65.1 423.45 ;
        RECT  63.9 433.05 65.1 434.85 ;
        RECT  59.1 433.95 60.3 434.85 ;
        RECT  59.1 421.05 60.3 422.25 ;
        RECT  61.5 423.3 62.7 432.75 ;
        RECT  57.3 428.1 59.4 429.0 ;
        RECT  62.7 428.1 66.9 429.0 ;
        RECT  59.1 429.15 60.3 430.35 ;
        RECT  61.5 429.15 62.7 430.35 ;
        RECT  59.1 428.25 60.3 429.45 ;
        RECT  61.5 428.25 62.7 429.45 ;
        RECT  63.9 423.45 65.1 424.65 ;
        RECT  63.9 433.95 65.1 435.15 ;
        RECT  59.4 429.15 60.6 430.35 ;
        RECT  66.9 434.85 78.9 435.75 ;
        RECT  66.9 420.15 78.9 421.05 ;
        RECT  75.9 420.6 76.8 423.45 ;
        RECT  75.9 432.9 76.8 435.3 ;
        RECT  68.85 420.6 69.75 423.45 ;
        RECT  73.65 420.6 74.55 423.45 ;
        RECT  68.85 432.45 69.75 435.3 ;
        RECT  66.9 425.7 69.0 426.6 ;
        RECT  66.9 429.0 72.0 429.9 ;
        RECT  74.55 428.1 78.9 429.0 ;
        RECT  68.7 427.65 69.9 428.85 ;
        RECT  71.1 427.65 72.3 428.85 ;
        RECT  71.1 427.65 72.3 428.85 ;
        RECT  73.5 427.65 74.7 428.85 ;
        RECT  68.7 428.25 69.9 429.45 ;
        RECT  71.1 428.25 72.3 429.45 ;
        RECT  71.1 428.25 72.3 429.45 ;
        RECT  73.5 428.25 74.7 429.45 ;
        RECT  75.9 423.45 77.1 424.65 ;
        RECT  75.9 433.65 77.1 434.85 ;
        RECT  74.1 440.7 75.0 441.6 ;
        RECT  71.1 440.7 72.0 441.6 ;
        RECT  74.1 433.65 75.0 441.15 ;
        RECT  71.55 440.7 74.55 441.6 ;
        RECT  71.1 441.15 72.0 443.85 ;
        RECT  69.0 426.9 70.2 428.1 ;
        RECT  72.0 430.2 73.2 431.4 ;
        RECT  78.9 434.85 88.5 435.75 ;
        RECT  78.9 420.15 88.5 421.05 ;
        RECT  85.5 421.05 86.7 423.45 ;
        RECT  85.5 433.05 86.7 434.85 ;
        RECT  80.7 433.95 81.9 434.85 ;
        RECT  80.7 421.05 81.9 422.25 ;
        RECT  83.1 423.3 84.3 432.75 ;
        RECT  78.9 428.1 81.0 429.0 ;
        RECT  84.3 428.1 88.5 429.0 ;
        RECT  80.7 429.15 81.9 430.35 ;
        RECT  83.1 429.15 84.3 430.35 ;
        RECT  80.7 428.25 81.9 429.45 ;
        RECT  83.1 428.25 84.3 429.45 ;
        RECT  85.5 423.45 86.7 424.65 ;
        RECT  85.5 433.95 86.7 435.15 ;
        RECT  81.0 429.15 82.2 430.35 ;
        RECT  66.9 425.4 68.1 426.6 ;
        RECT  51.0 425.4 52.2 426.6 ;
        RECT  17.25 39.0 18.15 79.8 ;
        RECT  71.7 39.0 72.6 79.8 ;
        RECT  71.7 69.0 72.6 80.4 ;
        RECT  68.4 79.2 71.7 80.4 ;
        RECT  69.9 71.4 70.8 78.0 ;
        RECT  69.6 75.0 69.9 78.0 ;
        RECT  69.6 71.4 69.9 72.6 ;
        RECT  67.2 76.2 68.4 80.4 ;
        RECT  67.2 69.0 68.4 72.6 ;
        RECT  63.6 79.2 67.2 80.4 ;
        RECT  66.3 73.8 67.2 75.0 ;
        RECT  66.0 72.6 66.3 75.0 ;
        RECT  65.1 71.4 66.0 78.0 ;
        RECT  64.8 76.2 65.1 78.0 ;
        RECT  64.8 71.4 65.1 72.6 ;
        RECT  62.4 76.2 63.6 80.4 ;
        RECT  48.6 79.2 62.4 80.4 ;
        RECT  61.8 73.5 64.2 74.7 ;
        RECT  63.6 69.0 67.2 69.9 ;
        RECT  62.4 69.0 63.6 72.6 ;
        RECT  61.2 69.0 62.4 70.2 ;
        RECT  58.8 76.8 60.0 78.0 ;
        RECT  59.7 73.5 60.9 75.9 ;
        RECT  57.9 71.4 58.8 78.0 ;
        RECT  57.6 76.2 57.9 78.0 ;
        RECT  57.6 71.4 57.9 72.6 ;
        RECT  55.5 71.4 56.4 78.0 ;
        RECT  55.2 76.2 55.5 78.0 ;
        RECT  55.2 71.4 55.5 73.8 ;
        RECT  53.1 71.4 54.0 78.0 ;
        RECT  52.8 76.2 53.1 78.0 ;
        RECT  52.8 71.4 53.1 73.8 ;
        RECT  51.0 73.8 51.9 75.0 ;
        RECT  50.1 71.4 51.0 78.0 ;
        RECT  49.8 75.0 50.1 78.0 ;
        RECT  49.8 71.4 50.1 72.6 ;
        RECT  47.4 76.2 48.6 80.4 ;
        RECT  42.9 79.2 47.4 80.4 ;
        RECT  46.5 74.1 48.9 75.3 ;
        RECT  48.6 69.0 61.2 69.9 ;
        RECT  47.4 69.0 48.6 72.6 ;
        RECT  45.3 76.8 46.5 78.0 ;
        RECT  44.4 71.4 45.3 78.0 ;
        RECT  44.1 76.2 44.4 78.0 ;
        RECT  44.1 71.4 44.4 72.6 ;
        RECT  42.9 69.0 47.4 69.9 ;
        RECT  41.7 76.2 42.9 80.4 ;
        RECT  38.1 79.2 41.7 80.4 ;
        RECT  40.8 73.5 42.0 74.7 ;
        RECT  41.7 69.0 42.9 72.6 ;
        RECT  40.5 72.6 40.8 78.0 ;
        RECT  39.9 71.4 40.5 78.0 ;
        RECT  39.3 76.2 39.9 78.0 ;
        RECT  39.6 71.4 39.9 73.8 ;
        RECT  39.3 71.4 39.6 72.6 ;
        RECT  36.9 76.2 38.1 80.4 ;
        RECT  21.9 79.2 36.9 80.4 ;
        RECT  36.3 73.5 38.7 74.7 ;
        RECT  38.1 69.0 41.7 69.9 ;
        RECT  36.9 69.0 38.1 72.6 ;
        RECT  35.7 69.0 36.9 70.2 ;
        RECT  32.4 76.8 33.6 78.0 ;
        RECT  33.3 73.5 34.5 75.9 ;
        RECT  31.5 71.4 32.4 78.0 ;
        RECT  31.2 76.2 31.5 78.0 ;
        RECT  31.2 71.4 31.5 72.6 ;
        RECT  29.1 71.4 30.0 78.0 ;
        RECT  28.8 76.2 29.1 78.0 ;
        RECT  28.8 71.4 29.1 73.8 ;
        RECT  26.7 71.4 27.6 78.0 ;
        RECT  26.4 76.2 26.7 78.0 ;
        RECT  26.4 71.4 26.7 73.8 ;
        RECT  24.6 73.8 25.5 75.0 ;
        RECT  23.7 71.4 24.6 78.0 ;
        RECT  23.4 75.0 23.7 78.0 ;
        RECT  23.4 71.4 23.7 72.6 ;
        RECT  22.2 69.0 35.7 69.9 ;
        RECT  21.9 76.2 22.2 78.0 ;
        RECT  21.0 76.2 21.9 80.4 ;
        RECT  21.3 69.0 22.2 72.6 ;
        RECT  21.0 71.4 21.3 72.6 ;
        RECT  19.5 76.2 21.0 77.4 ;
        RECT  18.6 74.1 19.5 75.3 ;
        RECT  17.7 69.0 18.6 80.4 ;
        RECT  71.7 58.8 72.6 70.2 ;
        RECT  68.4 58.8 71.7 60.0 ;
        RECT  69.9 61.2 70.8 67.8 ;
        RECT  69.6 61.2 69.9 64.2 ;
        RECT  69.6 66.6 69.9 67.8 ;
        RECT  67.2 58.8 68.4 63.0 ;
        RECT  67.2 66.6 68.4 70.2 ;
        RECT  63.6 58.8 67.2 60.0 ;
        RECT  66.3 64.2 67.2 65.4 ;
        RECT  66.0 64.2 66.3 66.6 ;
        RECT  65.1 61.2 66.0 67.8 ;
        RECT  64.8 61.2 65.1 63.0 ;
        RECT  64.8 66.6 65.1 67.8 ;
        RECT  62.4 58.8 63.6 63.0 ;
        RECT  48.6 58.8 62.4 60.0 ;
        RECT  61.8 64.5 64.2 65.7 ;
        RECT  63.6 69.3 67.2 70.2 ;
        RECT  62.4 66.6 63.6 70.2 ;
        RECT  61.2 69.0 62.4 70.2 ;
        RECT  58.8 61.2 60.0 62.4 ;
        RECT  59.7 63.3 60.9 65.7 ;
        RECT  57.9 61.2 58.8 67.8 ;
        RECT  57.6 61.2 57.9 63.0 ;
        RECT  57.6 66.6 57.9 67.8 ;
        RECT  55.5 61.2 56.4 67.8 ;
        RECT  55.2 61.2 55.5 63.0 ;
        RECT  55.2 65.4 55.5 67.8 ;
        RECT  53.1 61.2 54.0 67.8 ;
        RECT  52.8 61.2 53.1 63.0 ;
        RECT  52.8 65.4 53.1 67.8 ;
        RECT  51.0 64.2 51.9 65.4 ;
        RECT  50.1 61.2 51.0 67.8 ;
        RECT  49.8 61.2 50.1 64.2 ;
        RECT  49.8 66.6 50.1 67.8 ;
        RECT  47.4 58.8 48.6 63.0 ;
        RECT  42.9 58.8 47.4 60.0 ;
        RECT  46.5 63.9 48.9 65.1 ;
        RECT  48.6 69.3 61.2 70.2 ;
        RECT  47.4 66.6 48.6 70.2 ;
        RECT  45.3 61.2 46.5 62.4 ;
        RECT  44.4 61.2 45.3 67.8 ;
        RECT  44.1 61.2 44.4 63.0 ;
        RECT  44.1 66.6 44.4 67.8 ;
        RECT  42.9 69.3 47.4 70.2 ;
        RECT  41.7 58.8 42.9 63.0 ;
        RECT  38.1 58.8 41.7 60.0 ;
        RECT  40.8 64.5 42.0 65.7 ;
        RECT  41.7 66.6 42.9 70.2 ;
        RECT  40.5 61.2 40.8 66.6 ;
        RECT  39.9 61.2 40.5 67.8 ;
        RECT  39.3 61.2 39.9 63.0 ;
        RECT  39.6 65.4 39.9 67.8 ;
        RECT  39.3 66.6 39.6 67.8 ;
        RECT  36.9 58.8 38.1 63.0 ;
        RECT  21.9 58.8 36.9 60.0 ;
        RECT  36.3 64.5 38.7 65.7 ;
        RECT  38.1 69.3 41.7 70.2 ;
        RECT  36.9 66.6 38.1 70.2 ;
        RECT  35.7 69.0 36.9 70.2 ;
        RECT  32.4 61.2 33.6 62.4 ;
        RECT  33.3 63.3 34.5 65.7 ;
        RECT  31.5 61.2 32.4 67.8 ;
        RECT  31.2 61.2 31.5 63.0 ;
        RECT  31.2 66.6 31.5 67.8 ;
        RECT  29.1 61.2 30.0 67.8 ;
        RECT  28.8 61.2 29.1 63.0 ;
        RECT  28.8 65.4 29.1 67.8 ;
        RECT  26.7 61.2 27.6 67.8 ;
        RECT  26.4 61.2 26.7 63.0 ;
        RECT  26.4 65.4 26.7 67.8 ;
        RECT  24.6 64.2 25.5 65.4 ;
        RECT  23.7 61.2 24.6 67.8 ;
        RECT  23.4 61.2 23.7 64.2 ;
        RECT  23.4 66.6 23.7 67.8 ;
        RECT  22.2 69.3 35.7 70.2 ;
        RECT  21.9 61.2 22.2 63.0 ;
        RECT  21.0 58.8 21.9 63.0 ;
        RECT  21.3 66.6 22.2 70.2 ;
        RECT  21.0 66.6 21.3 67.8 ;
        RECT  19.5 61.8 21.0 63.0 ;
        RECT  18.6 63.9 19.5 65.1 ;
        RECT  17.7 58.8 18.6 70.2 ;
        RECT  71.7 48.6 72.6 60.0 ;
        RECT  68.4 58.8 71.7 60.0 ;
        RECT  69.9 51.0 70.8 57.6 ;
        RECT  69.6 54.6 69.9 57.6 ;
        RECT  69.6 51.0 69.9 52.2 ;
        RECT  67.2 55.8 68.4 60.0 ;
        RECT  67.2 48.6 68.4 52.2 ;
        RECT  63.6 58.8 67.2 60.0 ;
        RECT  66.3 53.4 67.2 54.6 ;
        RECT  66.0 52.2 66.3 54.6 ;
        RECT  65.1 51.0 66.0 57.6 ;
        RECT  64.8 55.8 65.1 57.6 ;
        RECT  64.8 51.0 65.1 52.2 ;
        RECT  62.4 55.8 63.6 60.0 ;
        RECT  48.6 58.8 62.4 60.0 ;
        RECT  61.8 53.1 64.2 54.3 ;
        RECT  63.6 48.6 67.2 49.5 ;
        RECT  62.4 48.6 63.6 52.2 ;
        RECT  61.2 48.6 62.4 49.8 ;
        RECT  58.8 56.4 60.0 57.6 ;
        RECT  59.7 53.1 60.9 55.5 ;
        RECT  57.9 51.0 58.8 57.6 ;
        RECT  57.6 55.8 57.9 57.6 ;
        RECT  57.6 51.0 57.9 52.2 ;
        RECT  55.5 51.0 56.4 57.6 ;
        RECT  55.2 55.8 55.5 57.6 ;
        RECT  55.2 51.0 55.5 53.4 ;
        RECT  53.1 51.0 54.0 57.6 ;
        RECT  52.8 55.8 53.1 57.6 ;
        RECT  52.8 51.0 53.1 53.4 ;
        RECT  51.0 53.4 51.9 54.6 ;
        RECT  50.1 51.0 51.0 57.6 ;
        RECT  49.8 54.6 50.1 57.6 ;
        RECT  49.8 51.0 50.1 52.2 ;
        RECT  47.4 55.8 48.6 60.0 ;
        RECT  42.9 58.8 47.4 60.0 ;
        RECT  46.5 53.7 48.9 54.9 ;
        RECT  48.6 48.6 61.2 49.5 ;
        RECT  47.4 48.6 48.6 52.2 ;
        RECT  45.3 56.4 46.5 57.6 ;
        RECT  44.4 51.0 45.3 57.6 ;
        RECT  44.1 55.8 44.4 57.6 ;
        RECT  44.1 51.0 44.4 52.2 ;
        RECT  42.9 48.6 47.4 49.5 ;
        RECT  41.7 55.8 42.9 60.0 ;
        RECT  38.1 58.8 41.7 60.0 ;
        RECT  40.8 53.1 42.0 54.3 ;
        RECT  41.7 48.6 42.9 52.2 ;
        RECT  40.5 52.2 40.8 57.6 ;
        RECT  39.9 51.0 40.5 57.6 ;
        RECT  39.3 55.8 39.9 57.6 ;
        RECT  39.6 51.0 39.9 53.4 ;
        RECT  39.3 51.0 39.6 52.2 ;
        RECT  36.9 55.8 38.1 60.0 ;
        RECT  21.9 58.8 36.9 60.0 ;
        RECT  36.3 53.1 38.7 54.3 ;
        RECT  38.1 48.6 41.7 49.5 ;
        RECT  36.9 48.6 38.1 52.2 ;
        RECT  35.7 48.6 36.9 49.8 ;
        RECT  32.4 56.4 33.6 57.6 ;
        RECT  33.3 53.1 34.5 55.5 ;
        RECT  31.5 51.0 32.4 57.6 ;
        RECT  31.2 55.8 31.5 57.6 ;
        RECT  31.2 51.0 31.5 52.2 ;
        RECT  29.1 51.0 30.0 57.6 ;
        RECT  28.8 55.8 29.1 57.6 ;
        RECT  28.8 51.0 29.1 53.4 ;
        RECT  26.7 51.0 27.6 57.6 ;
        RECT  26.4 55.8 26.7 57.6 ;
        RECT  26.4 51.0 26.7 53.4 ;
        RECT  24.6 53.4 25.5 54.6 ;
        RECT  23.7 51.0 24.6 57.6 ;
        RECT  23.4 54.6 23.7 57.6 ;
        RECT  23.4 51.0 23.7 52.2 ;
        RECT  22.2 48.6 35.7 49.5 ;
        RECT  21.9 55.8 22.2 57.6 ;
        RECT  21.0 55.8 21.9 60.0 ;
        RECT  21.3 48.6 22.2 52.2 ;
        RECT  21.0 51.0 21.3 52.2 ;
        RECT  19.5 55.8 21.0 57.0 ;
        RECT  18.6 53.7 19.5 54.9 ;
        RECT  17.7 48.6 18.6 60.0 ;
        RECT  71.7 38.4 72.6 49.8 ;
        RECT  68.4 38.4 71.7 39.6 ;
        RECT  69.9 40.8 70.8 47.4 ;
        RECT  69.6 40.8 69.9 43.8 ;
        RECT  69.6 46.2 69.9 47.4 ;
        RECT  67.2 38.4 68.4 42.6 ;
        RECT  67.2 46.2 68.4 49.8 ;
        RECT  63.6 38.4 67.2 39.6 ;
        RECT  66.3 43.8 67.2 45.0 ;
        RECT  66.0 43.8 66.3 46.2 ;
        RECT  65.1 40.8 66.0 47.4 ;
        RECT  64.8 40.8 65.1 42.6 ;
        RECT  64.8 46.2 65.1 47.4 ;
        RECT  62.4 38.4 63.6 42.6 ;
        RECT  48.6 38.4 62.4 39.6 ;
        RECT  61.8 44.1 64.2 45.3 ;
        RECT  63.6 48.9 67.2 49.8 ;
        RECT  62.4 46.2 63.6 49.8 ;
        RECT  61.2 48.6 62.4 49.8 ;
        RECT  58.8 40.8 60.0 42.0 ;
        RECT  59.7 42.9 60.9 45.3 ;
        RECT  57.9 40.8 58.8 47.4 ;
        RECT  57.6 40.8 57.9 42.6 ;
        RECT  57.6 46.2 57.9 47.4 ;
        RECT  55.5 40.8 56.4 47.4 ;
        RECT  55.2 40.8 55.5 42.6 ;
        RECT  55.2 45.0 55.5 47.4 ;
        RECT  53.1 40.8 54.0 47.4 ;
        RECT  52.8 40.8 53.1 42.6 ;
        RECT  52.8 45.0 53.1 47.4 ;
        RECT  51.0 43.8 51.9 45.0 ;
        RECT  50.1 40.8 51.0 47.4 ;
        RECT  49.8 40.8 50.1 43.8 ;
        RECT  49.8 46.2 50.1 47.4 ;
        RECT  47.4 38.4 48.6 42.6 ;
        RECT  42.9 38.4 47.4 39.6 ;
        RECT  46.5 43.5 48.9 44.7 ;
        RECT  48.6 48.9 61.2 49.8 ;
        RECT  47.4 46.2 48.6 49.8 ;
        RECT  45.3 40.8 46.5 42.0 ;
        RECT  44.4 40.8 45.3 47.4 ;
        RECT  44.1 40.8 44.4 42.6 ;
        RECT  44.1 46.2 44.4 47.4 ;
        RECT  42.9 48.9 47.4 49.8 ;
        RECT  41.7 38.4 42.9 42.6 ;
        RECT  38.1 38.4 41.7 39.6 ;
        RECT  40.8 44.1 42.0 45.3 ;
        RECT  41.7 46.2 42.9 49.8 ;
        RECT  40.5 40.8 40.8 46.2 ;
        RECT  39.9 40.8 40.5 47.4 ;
        RECT  39.3 40.8 39.9 42.6 ;
        RECT  39.6 45.0 39.9 47.4 ;
        RECT  39.3 46.2 39.6 47.4 ;
        RECT  36.9 38.4 38.1 42.6 ;
        RECT  21.9 38.4 36.9 39.6 ;
        RECT  36.3 44.1 38.7 45.3 ;
        RECT  38.1 48.9 41.7 49.8 ;
        RECT  36.9 46.2 38.1 49.8 ;
        RECT  35.7 48.6 36.9 49.8 ;
        RECT  32.4 40.8 33.6 42.0 ;
        RECT  33.3 42.9 34.5 45.3 ;
        RECT  31.5 40.8 32.4 47.4 ;
        RECT  31.2 40.8 31.5 42.6 ;
        RECT  31.2 46.2 31.5 47.4 ;
        RECT  29.1 40.8 30.0 47.4 ;
        RECT  28.8 40.8 29.1 42.6 ;
        RECT  28.8 45.0 29.1 47.4 ;
        RECT  26.7 40.8 27.6 47.4 ;
        RECT  26.4 40.8 26.7 42.6 ;
        RECT  26.4 45.0 26.7 47.4 ;
        RECT  24.6 43.8 25.5 45.0 ;
        RECT  23.7 40.8 24.6 47.4 ;
        RECT  23.4 40.8 23.7 43.8 ;
        RECT  23.4 46.2 23.7 47.4 ;
        RECT  22.2 48.9 35.7 49.8 ;
        RECT  21.9 40.8 22.2 42.6 ;
        RECT  21.0 38.4 21.9 42.6 ;
        RECT  21.3 46.2 22.2 49.8 ;
        RECT  21.0 46.2 21.3 47.4 ;
        RECT  19.5 41.4 21.0 42.6 ;
        RECT  18.6 43.5 19.5 44.7 ;
        RECT  17.7 38.4 18.6 49.8 ;
        RECT  88.5 202.35 89.4 203.25 ;
        RECT  88.95 202.35 124.35 203.25 ;
        RECT  88.5 202.8 89.4 208.2 ;
        RECT  88.5 226.35 89.4 227.25 ;
        RECT  88.95 226.35 124.35 227.25 ;
        RECT  88.5 221.4 89.4 226.8 ;
        RECT  88.5 231.75 89.4 232.65 ;
        RECT  88.95 231.75 124.35 232.65 ;
        RECT  88.5 232.2 89.4 237.6 ;
        RECT  88.5 255.75 89.4 256.65 ;
        RECT  88.95 255.75 124.35 256.65 ;
        RECT  88.5 250.8 89.4 256.2 ;
        RECT  88.5 261.15 89.4 262.05 ;
        RECT  88.95 261.15 124.35 262.05 ;
        RECT  88.5 261.6 89.4 267.0 ;
        RECT  88.5 285.15 89.4 286.05 ;
        RECT  88.95 285.15 124.35 286.05 ;
        RECT  88.5 280.2 89.4 285.6 ;
        RECT  88.5 290.55 89.4 291.45 ;
        RECT  88.95 290.55 124.35 291.45 ;
        RECT  88.5 291.0 89.4 296.4 ;
        RECT  88.5 314.55 89.4 315.45 ;
        RECT  88.95 314.55 124.35 315.45 ;
        RECT  88.5 309.6 89.4 315.0 ;
        RECT  88.5 319.95 89.4 320.85 ;
        RECT  88.95 319.95 124.35 320.85 ;
        RECT  88.5 320.4 89.4 325.8 ;
        RECT  88.5 343.95 89.4 344.85 ;
        RECT  88.95 343.95 124.35 344.85 ;
        RECT  88.5 339.0 89.4 344.4 ;
        RECT  88.5 349.35 89.4 350.25 ;
        RECT  88.95 349.35 124.35 350.25 ;
        RECT  88.5 349.8 89.4 355.2 ;
        RECT  88.5 373.35 89.4 374.25 ;
        RECT  88.95 373.35 124.35 374.25 ;
        RECT  88.5 368.4 89.4 373.8 ;
        RECT  88.5 378.75 89.4 379.65 ;
        RECT  88.95 378.75 124.35 379.65 ;
        RECT  88.5 379.2 89.4 384.6 ;
        RECT  88.5 402.75 89.4 403.65 ;
        RECT  88.95 402.75 124.35 403.65 ;
        RECT  88.5 397.8 89.4 403.2 ;
        RECT  88.5 408.15 89.4 409.05 ;
        RECT  88.95 408.15 124.35 409.05 ;
        RECT  88.5 408.6 89.4 414.0 ;
        RECT  88.5 432.15 89.4 433.05 ;
        RECT  88.95 432.15 124.35 433.05 ;
        RECT  88.5 427.2 89.4 432.6 ;
        RECT  90.6 88.8 91.8 90.0 ;
        RECT  87.9 104.7 89.1 105.9 ;
        RECT  85.2 147.6 86.4 148.8 ;
        RECT  82.5 163.5 83.7 164.7 ;
        RECT  114.0 33.3 115.2 34.5 ;
        RECT  108.6 28.65 109.8 29.85 ;
        RECT  111.3 26.25 112.5 27.45 ;
        RECT  114.0 446.4 115.2 447.6 ;
        RECT  116.7 97.95 117.9 99.15 ;
        RECT  119.4 196.05 120.6 197.25 ;
        RECT  16.5 76.5 17.7 77.7 ;
        RECT  53.7 456.6 54.6 457.5 ;
        RECT  53.7 435.3 54.6 457.05 ;
        RECT  54.15 456.6 107.25 457.5 ;
        RECT  105.9 456.6 107.1 457.8 ;
        RECT  71.7 35.85 72.6 36.75 ;
        RECT  0.0 35.85 72.15 36.75 ;
        RECT  71.7 36.3 72.6 39.0 ;
        RECT  95.1 437.1 97.5 438.3 ;
        RECT  133.8 437.1 135.0 438.3 ;
        RECT  144.0 437.1 145.2 438.3 ;
        RECT  154.2 437.1 155.4 438.3 ;
        RECT  122.7 437.1 123.9 438.3 ;
        RECT  101.7 8.1 104.1 9.3 ;
        RECT  133.5 8.1 134.7 9.3 ;
        RECT  133.5 8.1 134.7 9.3 ;
        RECT  153.9 8.1 155.1 9.3 ;
        RECT  87.75 229.05 88.95 230.25 ;
        RECT  87.75 258.45 88.95 259.65 ;
        RECT  87.75 287.85 88.95 289.05 ;
        RECT  87.75 317.25 88.95 318.45 ;
        RECT  87.75 346.65 88.95 347.85 ;
        RECT  87.75 376.05 88.95 377.25 ;
        RECT  87.75 405.45 88.95 406.65 ;
        RECT  87.75 434.85 88.95 436.05 ;
        RECT  95.1 140.55 97.5 141.75 ;
        RECT  95.1 199.35 97.5 200.55 ;
        RECT  75.0 69.15 76.2 70.35 ;
        RECT  95.1 69.15 97.5 70.35 ;
        RECT  75.0 69.15 76.2 70.35 ;
        RECT  95.1 69.15 97.5 70.35 ;
        RECT  75.0 48.75 76.2 49.95 ;
        RECT  95.1 48.75 97.5 49.95 ;
        RECT  75.0 48.75 76.2 49.95 ;
        RECT  95.1 48.75 97.5 49.95 ;
        RECT  -30.6 180.0 -28.95 180.9 ;
        RECT  -44.85 180.0 -43.2 180.9 ;
        RECT  -40.5 145.5 -39.6 151.8 ;
        RECT  -43.95 145.5 -43.05 154.5 ;
        RECT  -64.35 145.5 -63.45 157.2 ;
        RECT  -48.75 145.5 -47.85 159.9 ;
        RECT  -17.1 153.6 -16.2 164.4 ;
        RECT  -13.8 161.7 -12.9 164.4 ;
        RECT  -27.15 161.7 -26.25 164.4 ;
        RECT  -32.7 153.6 -31.8 164.4 ;
        RECT  -34.5 156.3 -33.6 164.4 ;
        RECT  -47.55 161.7 -46.65 164.4 ;
        RECT  -42.0 159.0 -41.1 164.4 ;
        RECT  -40.2 156.3 -39.3 164.4 ;
        RECT  -30.6 189.6 -29.7 215.1 ;
        RECT  -44.1 208.8 -43.2 212.4 ;
        RECT  -14.7 199.2 -13.8 217.8 ;
        RECT  -7.95 264.75 -3.0 265.65 ;
        RECT  -22.65 88.5 -21.75 223.5 ;
        RECT  -52.05 180.0 -51.15 220.5 ;
        RECT  -66.3 141.9 -21.75 142.8 ;
        RECT  -7.95 88.5 -7.05 233.4 ;
        RECT  -37.35 180.0 -36.45 230.4 ;
        RECT  -61.2 87.9 -27.15 88.8 ;
        RECT  -66.3 87.45 -35.7 88.35 ;
        RECT  -66.3 141.9 -35.7 142.8 ;
        RECT  -66.9 141.9 -55.5 142.8 ;
        RECT  -66.9 138.6 -65.7 141.9 ;
        RECT  -64.5 140.1 -57.9 141.0 ;
        RECT  -64.5 139.8 -61.5 140.1 ;
        RECT  -59.1 139.8 -57.9 140.1 ;
        RECT  -66.9 137.4 -62.7 138.6 ;
        RECT  -59.1 137.4 -55.5 138.6 ;
        RECT  -66.9 133.8 -65.7 137.4 ;
        RECT  -61.5 136.5 -60.3 137.4 ;
        RECT  -61.5 136.2 -59.1 136.5 ;
        RECT  -64.5 135.3 -57.9 136.2 ;
        RECT  -64.5 135.0 -62.7 135.3 ;
        RECT  -59.1 135.0 -57.9 135.3 ;
        RECT  -66.9 132.6 -62.7 133.8 ;
        RECT  -66.9 118.8 -65.7 132.6 ;
        RECT  -61.2 132.0 -60.0 134.4 ;
        RECT  -56.4 133.8 -55.5 137.4 ;
        RECT  -59.1 132.6 -55.5 133.8 ;
        RECT  -56.7 131.4 -55.5 132.6 ;
        RECT  -64.5 129.0 -63.3 130.2 ;
        RECT  -62.4 129.9 -60.0 131.1 ;
        RECT  -64.5 128.1 -57.9 129.0 ;
        RECT  -64.5 127.8 -62.7 128.1 ;
        RECT  -59.1 127.8 -57.9 128.1 ;
        RECT  -64.5 125.7 -57.9 126.6 ;
        RECT  -64.5 125.4 -62.7 125.7 ;
        RECT  -60.3 125.4 -57.9 125.7 ;
        RECT  -64.5 123.3 -57.9 124.2 ;
        RECT  -64.5 123.0 -62.7 123.3 ;
        RECT  -60.3 123.0 -57.9 123.3 ;
        RECT  -61.5 121.2 -60.3 122.1 ;
        RECT  -64.5 120.3 -57.9 121.2 ;
        RECT  -64.5 120.0 -61.5 120.3 ;
        RECT  -59.1 120.0 -57.9 120.3 ;
        RECT  -66.9 117.6 -62.7 118.8 ;
        RECT  -66.9 113.1 -65.7 117.6 ;
        RECT  -61.8 116.7 -60.6 119.1 ;
        RECT  -56.4 118.8 -55.5 131.4 ;
        RECT  -59.1 117.6 -55.5 118.8 ;
        RECT  -64.5 115.5 -63.3 116.7 ;
        RECT  -64.5 114.6 -57.9 115.5 ;
        RECT  -64.5 114.3 -62.7 114.6 ;
        RECT  -59.1 114.3 -57.9 114.6 ;
        RECT  -56.4 113.1 -55.5 117.6 ;
        RECT  -66.9 111.9 -62.7 113.1 ;
        RECT  -66.9 108.3 -65.7 111.9 ;
        RECT  -61.2 111.0 -60.0 112.2 ;
        RECT  -59.1 111.9 -55.5 113.1 ;
        RECT  -64.5 110.7 -59.1 111.0 ;
        RECT  -64.5 110.1 -57.9 110.7 ;
        RECT  -64.5 109.5 -62.7 110.1 ;
        RECT  -60.3 109.8 -57.9 110.1 ;
        RECT  -59.1 109.5 -57.9 109.8 ;
        RECT  -66.9 107.1 -62.7 108.3 ;
        RECT  -66.9 92.1 -65.7 107.1 ;
        RECT  -61.2 106.5 -60.0 108.9 ;
        RECT  -56.4 108.3 -55.5 111.9 ;
        RECT  -59.1 107.1 -55.5 108.3 ;
        RECT  -56.7 105.9 -55.5 107.1 ;
        RECT  -64.5 102.6 -63.3 103.8 ;
        RECT  -62.4 103.5 -60.0 104.7 ;
        RECT  -64.5 101.7 -57.9 102.6 ;
        RECT  -64.5 101.4 -62.7 101.7 ;
        RECT  -59.1 101.4 -57.9 101.7 ;
        RECT  -64.5 99.3 -57.9 100.2 ;
        RECT  -64.5 99.0 -62.7 99.3 ;
        RECT  -60.3 99.0 -57.9 99.3 ;
        RECT  -64.5 96.9 -57.9 97.8 ;
        RECT  -64.5 96.6 -62.7 96.9 ;
        RECT  -60.3 96.6 -57.9 96.9 ;
        RECT  -61.5 94.8 -60.3 95.7 ;
        RECT  -64.5 93.9 -57.9 94.8 ;
        RECT  -64.5 93.6 -61.5 93.9 ;
        RECT  -59.1 93.6 -57.9 93.9 ;
        RECT  -56.4 92.4 -55.5 105.9 ;
        RECT  -64.5 92.1 -62.7 92.4 ;
        RECT  -66.9 91.2 -62.7 92.1 ;
        RECT  -59.1 91.5 -55.5 92.4 ;
        RECT  -59.1 91.2 -57.9 91.5 ;
        RECT  -63.9 89.7 -62.7 91.2 ;
        RECT  -61.8 88.8 -60.6 89.7 ;
        RECT  -66.9 87.9 -55.5 88.8 ;
        RECT  -56.7 141.9 -45.3 142.8 ;
        RECT  -46.5 138.6 -45.3 141.9 ;
        RECT  -54.3 140.1 -47.7 141.0 ;
        RECT  -50.7 139.8 -47.7 140.1 ;
        RECT  -54.3 139.8 -53.1 140.1 ;
        RECT  -49.5 137.4 -45.3 138.6 ;
        RECT  -56.7 137.4 -53.1 138.6 ;
        RECT  -46.5 133.8 -45.3 137.4 ;
        RECT  -51.9 136.5 -50.7 137.4 ;
        RECT  -53.1 136.2 -50.7 136.5 ;
        RECT  -54.3 135.3 -47.7 136.2 ;
        RECT  -49.5 135.0 -47.7 135.3 ;
        RECT  -54.3 135.0 -53.1 135.3 ;
        RECT  -49.5 132.6 -45.3 133.8 ;
        RECT  -46.5 118.8 -45.3 132.6 ;
        RECT  -52.2 132.0 -51.0 134.4 ;
        RECT  -56.7 133.8 -55.8 137.4 ;
        RECT  -56.7 132.6 -53.1 133.8 ;
        RECT  -56.7 131.4 -55.5 132.6 ;
        RECT  -48.9 129.0 -47.7 130.2 ;
        RECT  -52.2 129.9 -49.8 131.1 ;
        RECT  -54.3 128.1 -47.7 129.0 ;
        RECT  -49.5 127.8 -47.7 128.1 ;
        RECT  -54.3 127.8 -53.1 128.1 ;
        RECT  -54.3 125.7 -47.7 126.6 ;
        RECT  -49.5 125.4 -47.7 125.7 ;
        RECT  -54.3 125.4 -51.9 125.7 ;
        RECT  -54.3 123.3 -47.7 124.2 ;
        RECT  -49.5 123.0 -47.7 123.3 ;
        RECT  -54.3 123.0 -51.9 123.3 ;
        RECT  -51.9 121.2 -50.7 122.1 ;
        RECT  -54.3 120.3 -47.7 121.2 ;
        RECT  -50.7 120.0 -47.7 120.3 ;
        RECT  -54.3 120.0 -53.1 120.3 ;
        RECT  -49.5 117.6 -45.3 118.8 ;
        RECT  -46.5 113.1 -45.3 117.6 ;
        RECT  -51.6 116.7 -50.4 119.1 ;
        RECT  -56.7 118.8 -55.8 131.4 ;
        RECT  -56.7 117.6 -53.1 118.8 ;
        RECT  -48.9 115.5 -47.7 116.7 ;
        RECT  -54.3 114.6 -47.7 115.5 ;
        RECT  -49.5 114.3 -47.7 114.6 ;
        RECT  -54.3 114.3 -53.1 114.6 ;
        RECT  -56.7 113.1 -55.8 117.6 ;
        RECT  -49.5 111.9 -45.3 113.1 ;
        RECT  -46.5 108.3 -45.3 111.9 ;
        RECT  -52.2 111.0 -51.0 112.2 ;
        RECT  -56.7 111.9 -53.1 113.1 ;
        RECT  -53.1 110.7 -47.7 111.0 ;
        RECT  -54.3 110.1 -47.7 110.7 ;
        RECT  -49.5 109.5 -47.7 110.1 ;
        RECT  -54.3 109.8 -51.9 110.1 ;
        RECT  -54.3 109.5 -53.1 109.8 ;
        RECT  -49.5 107.1 -45.3 108.3 ;
        RECT  -46.5 92.1 -45.3 107.1 ;
        RECT  -52.2 106.5 -51.0 108.9 ;
        RECT  -56.7 108.3 -55.8 111.9 ;
        RECT  -56.7 107.1 -53.1 108.3 ;
        RECT  -56.7 105.9 -55.5 107.1 ;
        RECT  -48.9 102.6 -47.7 103.8 ;
        RECT  -52.2 103.5 -49.8 104.7 ;
        RECT  -54.3 101.7 -47.7 102.6 ;
        RECT  -49.5 101.4 -47.7 101.7 ;
        RECT  -54.3 101.4 -53.1 101.7 ;
        RECT  -54.3 99.3 -47.7 100.2 ;
        RECT  -49.5 99.0 -47.7 99.3 ;
        RECT  -54.3 99.0 -51.9 99.3 ;
        RECT  -54.3 96.9 -47.7 97.8 ;
        RECT  -49.5 96.6 -47.7 96.9 ;
        RECT  -54.3 96.6 -51.9 96.9 ;
        RECT  -51.9 94.8 -50.7 95.7 ;
        RECT  -54.3 93.9 -47.7 94.8 ;
        RECT  -50.7 93.6 -47.7 93.9 ;
        RECT  -54.3 93.6 -53.1 93.9 ;
        RECT  -56.7 92.4 -55.8 105.9 ;
        RECT  -49.5 92.1 -47.7 92.4 ;
        RECT  -49.5 91.2 -45.3 92.1 ;
        RECT  -56.7 91.5 -53.1 92.4 ;
        RECT  -54.3 91.2 -53.1 91.5 ;
        RECT  -49.5 89.7 -48.3 91.2 ;
        RECT  -51.6 88.8 -50.4 89.7 ;
        RECT  -56.7 87.9 -45.3 88.8 ;
        RECT  -46.5 141.9 -35.1 142.8 ;
        RECT  -46.5 138.6 -45.3 141.9 ;
        RECT  -44.1 140.1 -37.5 141.0 ;
        RECT  -44.1 139.8 -41.1 140.1 ;
        RECT  -38.7 139.8 -37.5 140.1 ;
        RECT  -46.5 137.4 -42.3 138.6 ;
        RECT  -38.7 137.4 -35.1 138.6 ;
        RECT  -46.5 133.8 -45.3 137.4 ;
        RECT  -41.1 136.5 -39.9 137.4 ;
        RECT  -41.1 136.2 -38.7 136.5 ;
        RECT  -44.1 135.3 -37.5 136.2 ;
        RECT  -44.1 135.0 -42.3 135.3 ;
        RECT  -38.7 135.0 -37.5 135.3 ;
        RECT  -46.5 132.6 -42.3 133.8 ;
        RECT  -46.5 118.8 -45.3 132.6 ;
        RECT  -40.8 132.0 -39.6 134.4 ;
        RECT  -36.0 133.8 -35.1 137.4 ;
        RECT  -38.7 132.6 -35.1 133.8 ;
        RECT  -36.3 131.4 -35.1 132.6 ;
        RECT  -44.1 129.0 -42.9 130.2 ;
        RECT  -42.0 129.9 -39.6 131.1 ;
        RECT  -44.1 128.1 -37.5 129.0 ;
        RECT  -44.1 127.8 -42.3 128.1 ;
        RECT  -38.7 127.8 -37.5 128.1 ;
        RECT  -44.1 125.7 -37.5 126.6 ;
        RECT  -44.1 125.4 -42.3 125.7 ;
        RECT  -39.9 125.4 -37.5 125.7 ;
        RECT  -44.1 123.3 -37.5 124.2 ;
        RECT  -44.1 123.0 -42.3 123.3 ;
        RECT  -39.9 123.0 -37.5 123.3 ;
        RECT  -41.1 121.2 -39.9 122.1 ;
        RECT  -44.1 120.3 -37.5 121.2 ;
        RECT  -44.1 120.0 -41.1 120.3 ;
        RECT  -38.7 120.0 -37.5 120.3 ;
        RECT  -46.5 117.6 -42.3 118.8 ;
        RECT  -46.5 113.1 -45.3 117.6 ;
        RECT  -41.4 116.7 -40.2 119.1 ;
        RECT  -36.0 118.8 -35.1 131.4 ;
        RECT  -38.7 117.6 -35.1 118.8 ;
        RECT  -44.1 115.5 -42.9 116.7 ;
        RECT  -44.1 114.6 -37.5 115.5 ;
        RECT  -44.1 114.3 -42.3 114.6 ;
        RECT  -38.7 114.3 -37.5 114.6 ;
        RECT  -36.0 113.1 -35.1 117.6 ;
        RECT  -46.5 111.9 -42.3 113.1 ;
        RECT  -46.5 108.3 -45.3 111.9 ;
        RECT  -40.8 111.0 -39.6 112.2 ;
        RECT  -38.7 111.9 -35.1 113.1 ;
        RECT  -44.1 110.7 -38.7 111.0 ;
        RECT  -44.1 110.1 -37.5 110.7 ;
        RECT  -44.1 109.5 -42.3 110.1 ;
        RECT  -39.9 109.8 -37.5 110.1 ;
        RECT  -38.7 109.5 -37.5 109.8 ;
        RECT  -46.5 107.1 -42.3 108.3 ;
        RECT  -46.5 92.1 -45.3 107.1 ;
        RECT  -40.8 106.5 -39.6 108.9 ;
        RECT  -36.0 108.3 -35.1 111.9 ;
        RECT  -38.7 107.1 -35.1 108.3 ;
        RECT  -36.3 105.9 -35.1 107.1 ;
        RECT  -44.1 102.6 -42.9 103.8 ;
        RECT  -42.0 103.5 -39.6 104.7 ;
        RECT  -44.1 101.7 -37.5 102.6 ;
        RECT  -44.1 101.4 -42.3 101.7 ;
        RECT  -38.7 101.4 -37.5 101.7 ;
        RECT  -44.1 99.3 -37.5 100.2 ;
        RECT  -44.1 99.0 -42.3 99.3 ;
        RECT  -39.9 99.0 -37.5 99.3 ;
        RECT  -44.1 96.9 -37.5 97.8 ;
        RECT  -44.1 96.6 -42.3 96.9 ;
        RECT  -39.9 96.6 -37.5 96.9 ;
        RECT  -41.1 94.8 -39.9 95.7 ;
        RECT  -44.1 93.9 -37.5 94.8 ;
        RECT  -44.1 93.6 -41.1 93.9 ;
        RECT  -38.7 93.6 -37.5 93.9 ;
        RECT  -36.0 92.4 -35.1 105.9 ;
        RECT  -44.1 92.1 -42.3 92.4 ;
        RECT  -46.5 91.2 -42.3 92.1 ;
        RECT  -38.7 91.5 -35.1 92.4 ;
        RECT  -38.7 91.2 -37.5 91.5 ;
        RECT  -43.5 89.7 -42.3 91.2 ;
        RECT  -41.4 88.8 -40.2 89.7 ;
        RECT  -46.5 87.9 -35.1 88.8 ;
        RECT  -7.95 128.7 -7.05 145.5 ;
        RECT  -22.65 128.7 -21.75 145.5 ;
        RECT  -21.75 142.5 -19.35 143.7 ;
        RECT  -9.75 142.5 -7.95 143.7 ;
        RECT  -19.5 132.9 -10.05 134.1 ;
        RECT  -19.5 137.7 -10.05 138.9 ;
        RECT  -14.7 128.7 -13.8 130.8 ;
        RECT  -14.7 138.9 -13.8 145.5 ;
        RECT  -11.25 130.5 -10.05 131.7 ;
        RECT  -11.25 132.9 -10.05 134.1 ;
        RECT  -11.25 135.3 -10.05 136.5 ;
        RECT  -11.25 137.7 -10.05 138.9 ;
        RECT  -11.25 140.1 -10.05 141.3 ;
        RECT  -13.05 130.5 -12.15 131.4 ;
        RECT  -13.05 135.3 -12.15 136.2 ;
        RECT  -13.05 135.3 -12.15 136.2 ;
        RECT  -13.05 140.1 -12.15 141.0 ;
        RECT  -12.15 130.5 -10.05 131.4 ;
        RECT  -12.6 130.5 -12.15 131.4 ;
        RECT  -13.05 130.95 -12.15 135.75 ;
        RECT  -12.6 135.3 -10.05 136.2 ;
        RECT  -12.15 135.3 -10.05 136.2 ;
        RECT  -12.6 135.3 -12.15 136.2 ;
        RECT  -13.05 135.75 -12.15 140.55 ;
        RECT  -12.6 140.1 -10.05 141.0 ;
        RECT  -9.15 132.9 -8.25 133.8 ;
        RECT  -9.15 137.7 -8.25 138.6 ;
        RECT  -10.05 132.9 -9.15 133.8 ;
        RECT  -9.15 132.9 -8.7 133.8 ;
        RECT  -9.15 133.35 -8.25 138.15 ;
        RECT  -10.05 137.7 -8.7 138.6 ;
        RECT  -20.55 130.5 -19.35 131.7 ;
        RECT  -20.55 132.9 -19.35 134.1 ;
        RECT  -20.55 135.3 -19.35 136.5 ;
        RECT  -20.55 137.7 -19.35 138.9 ;
        RECT  -20.55 140.1 -19.35 141.3 ;
        RECT  -22.35 130.5 -21.45 131.4 ;
        RECT  -22.35 135.3 -21.45 136.2 ;
        RECT  -22.35 135.3 -21.45 136.2 ;
        RECT  -22.35 140.1 -21.45 141.0 ;
        RECT  -21.45 130.5 -19.35 131.4 ;
        RECT  -21.9 130.5 -21.45 131.4 ;
        RECT  -22.35 130.95 -21.45 135.75 ;
        RECT  -21.9 135.3 -19.35 136.2 ;
        RECT  -21.45 135.3 -19.35 136.2 ;
        RECT  -21.9 135.3 -21.45 136.2 ;
        RECT  -22.35 135.75 -21.45 140.55 ;
        RECT  -21.9 140.1 -19.35 141.0 ;
        RECT  -18.45 132.9 -17.55 133.8 ;
        RECT  -18.45 137.7 -17.55 138.6 ;
        RECT  -19.35 132.9 -18.45 133.8 ;
        RECT  -18.45 132.9 -18.0 133.8 ;
        RECT  -18.45 133.35 -17.55 138.15 ;
        RECT  -19.35 137.7 -18.0 138.6 ;
        RECT  -20.55 142.5 -19.35 143.7 ;
        RECT  -10.05 142.5 -8.85 143.7 ;
        RECT  -14.85 130.8 -13.65 132.0 ;
        RECT  -7.95 88.5 -7.05 119.7 ;
        RECT  -22.65 88.5 -21.75 119.7 ;
        RECT  -14.1 116.4 -13.2 119.7 ;
        RECT  -16.05 102.0 -15.15 119.7 ;
        RECT  -22.2 90.6 -19.65 91.5 ;
        RECT  -8.85 109.8 -7.5 110.7 ;
        RECT  -21.75 117.0 -19.65 117.9 ;
        RECT  -21.75 112.2 -19.65 113.1 ;
        RECT  -21.75 107.4 -19.65 108.3 ;
        RECT  -8.85 117.0 -7.05 117.9 ;
        RECT  -8.85 112.2 -7.05 113.1 ;
        RECT  -13.65 116.7 -12.45 117.9 ;
        RECT  -13.65 114.3 -12.45 115.5 ;
        RECT  -13.65 114.3 -12.45 115.5 ;
        RECT  -13.65 111.9 -12.45 113.1 ;
        RECT  -16.05 116.7 -14.85 117.9 ;
        RECT  -16.05 114.3 -14.85 115.5 ;
        RECT  -16.05 111.9 -14.85 113.1 ;
        RECT  -16.05 109.5 -14.85 110.7 ;
        RECT  -16.05 107.1 -14.85 108.3 ;
        RECT  -16.05 102.3 -14.85 103.5 ;
        RECT  -16.05 99.9 -14.85 101.1 ;
        RECT  -16.05 97.5 -14.85 98.7 ;
        RECT  -16.05 95.1 -14.85 96.3 ;
        RECT  -16.05 92.7 -14.85 93.9 ;
        RECT  -19.65 90.3 -18.45 91.5 ;
        RECT  -8.85 109.5 -7.65 110.7 ;
        RECT  -13.05 116.4 -11.85 117.6 ;
        RECT  -15.0 102.0 -13.8 103.2 ;
        RECT  -14.1 114.45 -13.2 115.35 ;
        RECT  -14.1 88.5 -13.2 114.9 ;
        RECT  -18.45 114.45 -13.65 115.35 ;
        RECT  -19.65 99.9 -18.45 101.1 ;
        RECT  -14.1 100.05 -13.2 100.95 ;
        RECT  -14.1 88.5 -13.2 100.5 ;
        RECT  -14.25 99.9 -13.05 101.1 ;
        RECT  -19.65 95.1 -18.45 96.3 ;
        RECT  -14.1 95.25 -13.2 96.15 ;
        RECT  -14.1 88.5 -13.2 95.7 ;
        RECT  -14.25 95.1 -13.05 96.3 ;
        RECT  -22.2 114.45 -21.3 115.35 ;
        RECT  -21.75 114.45 -19.65 115.35 ;
        RECT  -22.2 105.3 -21.3 114.9 ;
        RECT  -22.2 109.65 -21.3 110.55 ;
        RECT  -21.75 109.65 -19.65 110.55 ;
        RECT  -22.2 105.3 -21.3 110.1 ;
        RECT  -22.2 102.45 -21.3 103.35 ;
        RECT  -21.75 102.45 -19.65 103.35 ;
        RECT  -22.2 102.9 -21.3 105.3 ;
        RECT  -22.2 97.65 -21.3 98.55 ;
        RECT  -21.75 97.65 -19.65 98.55 ;
        RECT  -22.2 98.1 -21.3 105.3 ;
        RECT  -22.2 92.85 -21.3 93.75 ;
        RECT  -21.75 92.85 -19.65 93.75 ;
        RECT  -22.2 93.3 -21.3 105.3 ;
        RECT  -7.95 164.4 -7.05 176.4 ;
        RECT  -22.65 164.4 -21.75 176.4 ;
        RECT  -22.2 173.4 -19.35 174.3 ;
        RECT  -9.9 173.4 -7.5 174.3 ;
        RECT  -22.2 166.35 -19.35 167.25 ;
        RECT  -22.2 171.15 -19.35 172.05 ;
        RECT  -10.35 166.35 -7.5 167.25 ;
        RECT  -17.1 164.4 -16.2 166.5 ;
        RECT  -13.8 164.4 -12.9 169.5 ;
        RECT  -14.7 172.05 -13.8 176.4 ;
        RECT  -11.55 166.2 -10.35 167.4 ;
        RECT  -11.55 168.6 -10.35 169.8 ;
        RECT  -11.55 168.6 -10.35 169.8 ;
        RECT  -11.55 171.0 -10.35 172.2 ;
        RECT  -20.55 166.2 -19.35 167.4 ;
        RECT  -20.55 168.6 -19.35 169.8 ;
        RECT  -20.55 168.6 -19.35 169.8 ;
        RECT  -20.55 171.0 -19.35 172.2 ;
        RECT  -20.55 173.4 -19.35 174.6 ;
        RECT  -10.35 173.4 -9.15 174.6 ;
        RECT  -17.1 171.6 -16.2 172.5 ;
        RECT  -17.1 168.6 -16.2 169.5 ;
        RECT  -16.65 171.6 -9.15 172.5 ;
        RECT  -17.1 169.05 -16.2 172.05 ;
        RECT  -19.35 168.6 -16.65 169.5 ;
        RECT  -17.1 166.5 -15.9 167.7 ;
        RECT  -13.8 169.5 -12.6 170.7 ;
        RECT  -43.05 236.1 -41.85 237.3 ;
        RECT  -45.0 236.1 -44.1 237.0 ;
        RECT  -51.75 250.95 -49.2 251.85 ;
        RECT  -61.95 292.65 -7.95 293.55 ;
        RECT  -8.4 268.8 -7.5 288.0 ;
        RECT  -37.8 268.8 -36.9 288.0 ;
        RECT  -41.85 229.95 -32.25 230.85 ;
        RECT  -41.85 215.25 -32.25 216.15 ;
        RECT  -40.05 216.15 -38.85 219.9 ;
        RECT  -40.05 228.15 -38.85 229.95 ;
        RECT  -35.25 229.05 -34.05 229.95 ;
        RECT  -35.25 216.15 -34.05 217.2 ;
        RECT  -37.65 219.75 -36.45 227.85 ;
        RECT  -34.35 223.8 -32.25 224.7 ;
        RECT  -41.85 223.8 -37.65 224.7 ;
        RECT  -35.25 226.65 -34.05 227.85 ;
        RECT  -37.65 226.65 -36.45 227.85 ;
        RECT  -35.25 217.2 -34.05 219.9 ;
        RECT  -37.65 217.2 -36.45 219.9 ;
        RECT  -40.05 217.2 -38.85 219.9 ;
        RECT  -40.05 227.85 -38.85 229.05 ;
        RECT  -35.55 223.65 -34.35 224.85 ;
        RECT  -16.35 234.75 -15.15 235.95 ;
        RECT  -16.35 232.35 -15.15 233.55 ;
        RECT  -14.85 265.8 -13.65 267.0 ;
        RECT  -8.4 257.4 -7.5 267.0 ;
        RECT  -23.1 257.4 -22.2 267.0 ;
        RECT  -22.2 259.2 -18.45 260.4 ;
        RECT  -10.2 259.2 -8.4 260.4 ;
        RECT  -9.3 264.0 -8.4 265.2 ;
        RECT  -22.2 264.0 -21.15 265.2 ;
        RECT  -18.6 261.6 -10.5 262.8 ;
        RECT  -14.55 264.9 -13.65 267.0 ;
        RECT  -14.1 264.0 -12.9 265.2 ;
        RECT  -14.1 261.6 -12.9 262.8 ;
        RECT  -13.95 264.0 -11.25 265.2 ;
        RECT  -13.95 261.6 -11.25 262.8 ;
        RECT  -18.45 259.2 -15.75 260.4 ;
        RECT  -9.3 259.2 -8.1 260.4 ;
        RECT  -13.5 263.7 -12.3 264.9 ;
        RECT  -14.85 256.2 -13.65 257.4 ;
        RECT  -8.4 247.8 -7.5 257.4 ;
        RECT  -23.1 247.8 -22.2 257.4 ;
        RECT  -22.2 249.6 -18.45 250.8 ;
        RECT  -10.2 249.6 -8.4 250.8 ;
        RECT  -9.3 254.4 -8.4 255.6 ;
        RECT  -22.2 254.4 -21.15 255.6 ;
        RECT  -18.6 252.0 -10.5 253.2 ;
        RECT  -14.55 255.3 -13.65 257.4 ;
        RECT  -14.1 254.4 -12.9 255.6 ;
        RECT  -14.1 252.0 -12.9 253.2 ;
        RECT  -13.95 254.4 -11.25 255.6 ;
        RECT  -13.95 252.0 -11.25 253.2 ;
        RECT  -18.45 249.6 -15.75 250.8 ;
        RECT  -9.3 249.6 -8.1 250.8 ;
        RECT  -13.5 254.1 -12.3 255.3 ;
        RECT  -31.65 247.8 -30.45 249.0 ;
        RECT  -37.8 247.8 -36.9 257.4 ;
        RECT  -23.1 247.8 -22.2 257.4 ;
        RECT  -26.85 254.4 -23.1 255.6 ;
        RECT  -36.9 254.4 -35.1 255.6 ;
        RECT  -36.9 249.6 -36.0 250.8 ;
        RECT  -24.15 249.6 -23.1 250.8 ;
        RECT  -34.8 252.0 -26.7 253.2 ;
        RECT  -31.65 247.8 -30.75 249.9 ;
        RECT  -32.4 249.6 -31.2 250.8 ;
        RECT  -32.4 252.0 -31.2 253.2 ;
        RECT  -34.05 249.6 -31.35 250.8 ;
        RECT  -34.05 252.0 -31.35 253.2 ;
        RECT  -29.55 254.4 -26.85 255.6 ;
        RECT  -37.2 254.4 -36.0 255.6 ;
        RECT  -33.0 249.9 -31.8 251.1 ;
        RECT  -31.65 257.4 -30.45 258.6 ;
        RECT  -37.8 257.4 -36.9 267.0 ;
        RECT  -23.1 257.4 -22.2 267.0 ;
        RECT  -26.85 264.0 -23.1 265.2 ;
        RECT  -36.9 264.0 -35.1 265.2 ;
        RECT  -36.9 259.2 -36.0 260.4 ;
        RECT  -24.15 259.2 -23.1 260.4 ;
        RECT  -34.8 261.6 -26.7 262.8 ;
        RECT  -31.65 257.4 -30.75 259.5 ;
        RECT  -32.4 259.2 -31.2 260.4 ;
        RECT  -32.4 261.6 -31.2 262.8 ;
        RECT  -34.05 259.2 -31.35 260.4 ;
        RECT  -34.05 261.6 -31.35 262.8 ;
        RECT  -29.55 264.0 -26.85 265.2 ;
        RECT  -37.2 264.0 -36.0 265.2 ;
        RECT  -33.0 259.5 -31.8 260.7 ;
        RECT  -14.85 260.4 -13.65 261.6 ;
        RECT  -14.85 250.8 -13.65 252.0 ;
        RECT  -31.65 253.2 -30.45 254.4 ;
        RECT  -62.55 267.6 -51.75 268.8 ;
        RECT  -53.55 265.5 -52.35 267.6 ;
        RECT  -56.55 265.5 -55.35 266.7 ;
        RECT  -59.55 265.5 -58.35 266.7 ;
        RECT  -62.55 265.5 -61.35 267.6 ;
        RECT  -56.25 264.6 -55.05 265.5 ;
        RECT  -57.45 263.4 -52.35 264.6 ;
        RECT  -53.55 258.3 -52.35 263.4 ;
        RECT  -56.25 260.1 -55.05 263.4 ;
        RECT  -59.85 261.9 -58.65 265.5 ;
        RECT  -59.85 260.7 -58.05 261.9 ;
        RECT  -59.85 260.1 -58.65 260.7 ;
        RECT  -55.95 258.9 -54.75 260.1 ;
        RECT  -60.15 258.9 -58.95 260.1 ;
        RECT  -62.55 258.9 -61.35 264.6 ;
        RECT  -58.05 257.4 -56.85 257.7 ;
        RECT  -62.55 256.2 -51.75 257.4 ;
        RECT  -55.95 254.1 -53.25 255.3 ;
        RECT  -60.15 254.1 -57.45 255.3 ;
        RECT  -62.55 239.4 -51.15 240.6 ;
        RECT  -53.55 240.6 -52.35 242.7 ;
        RECT  -56.55 241.5 -55.35 242.7 ;
        RECT  -59.55 241.5 -58.35 242.7 ;
        RECT  -62.55 240.6 -61.35 242.7 ;
        RECT  -56.25 242.7 -55.05 243.6 ;
        RECT  -53.55 243.6 -52.35 249.3 ;
        RECT  -57.45 243.6 -55.05 244.8 ;
        RECT  -56.25 244.8 -55.05 248.1 ;
        RECT  -59.85 242.7 -58.65 246.3 ;
        RECT  -59.85 246.3 -58.05 247.5 ;
        RECT  -59.85 247.5 -58.65 248.1 ;
        RECT  -55.95 248.1 -54.75 249.3 ;
        RECT  -60.15 248.1 -58.95 249.3 ;
        RECT  -62.55 243.6 -61.35 249.3 ;
        RECT  -58.05 250.5 -56.85 250.8 ;
        RECT  -62.55 250.8 -51.15 252.0 ;
        RECT  -55.95 252.9 -53.25 254.1 ;
        RECT  -60.15 252.9 -57.45 254.1 ;
        RECT  -62.55 238.2 -51.15 239.4 ;
        RECT  -53.55 236.1 -52.35 238.2 ;
        RECT  -56.55 236.1 -55.35 237.3 ;
        RECT  -59.55 236.1 -58.35 237.3 ;
        RECT  -62.55 236.1 -61.35 238.2 ;
        RECT  -56.25 235.2 -55.05 236.1 ;
        RECT  -53.55 229.5 -52.35 235.2 ;
        RECT  -57.45 234.0 -55.05 235.2 ;
        RECT  -56.25 230.7 -55.05 234.0 ;
        RECT  -59.85 232.5 -58.65 236.1 ;
        RECT  -59.85 231.3 -58.05 232.5 ;
        RECT  -59.85 230.7 -58.65 231.3 ;
        RECT  -55.95 229.5 -54.75 230.7 ;
        RECT  -60.15 229.5 -58.95 230.7 ;
        RECT  -62.55 229.5 -61.35 235.2 ;
        RECT  -58.05 228.0 -56.85 228.3 ;
        RECT  -62.55 226.8 -51.15 228.0 ;
        RECT  -55.95 224.7 -53.25 225.9 ;
        RECT  -60.15 224.7 -57.45 225.9 ;
        RECT  -43.05 235.35 -41.85 236.55 ;
        RECT  -14.55 264.75 -13.65 265.65 ;
        RECT  -14.1 264.75 -7.95 265.65 ;
        RECT  -14.55 263.4 -13.65 265.2 ;
        RECT  -32.7 238.05 -31.8 238.95 ;
        RECT  -45.0 238.2 -44.1 239.1 ;
        RECT  -32.7 236.55 -31.8 238.65 ;
        RECT  -45.0 236.55 -44.1 238.65 ;
        RECT  -32.85 237.9 -31.65 239.1 ;
        RECT  -45.15 238.05 -43.95 239.25 ;
        RECT  -55.8 271.05 -54.9 271.95 ;
        RECT  -55.35 271.2 -44.55 272.1 ;
        RECT  -55.95 270.9 -54.75 272.1 ;
        RECT  -13.95 239.55 -12.75 240.75 ;
        RECT  -13.65 220.5 -12.75 221.4 ;
        RECT  -32.1 220.65 -31.2 221.55 ;
        RECT  -31.65 220.65 -13.2 221.55 ;
        RECT  -13.8 220.35 -12.6 221.55 ;
        RECT  -32.25 220.5 -31.05 221.7 ;
        RECT  -32.85 271.2 -31.65 272.4 ;
        RECT  -13.8 239.55 -12.6 240.75 ;
        RECT  -50.25 249.6 -49.05 250.8 ;
        RECT  -16.35 239.55 -15.45 240.45 ;
        RECT  -16.35 240.0 -15.45 242.55 ;
        RECT  -32.25 239.55 -15.9 240.45 ;
        RECT  -45.9 244.65 -45.0 245.55 ;
        RECT  -45.45 244.65 -32.25 245.55 ;
        RECT  -46.05 244.5 -44.85 245.7 ;
        RECT  -16.35 243.3 -15.45 244.2 ;
        RECT  -16.35 240.15 -15.45 243.75 ;
        RECT  -32.25 243.3 -15.9 244.2 ;
        RECT  -23.1 268.35 -22.2 269.25 ;
        RECT  -23.1 267.0 -22.2 268.8 ;
        RECT  -45.45 268.35 -22.65 269.25 ;
        RECT  -45.9 264.75 -45.0 265.65 ;
        RECT  -45.45 264.75 -22.65 265.65 ;
        RECT  -46.05 264.6 -44.85 265.8 ;
        RECT  -8.4 229.95 -7.5 230.85 ;
        RECT  -8.4 172.2 -7.5 173.1 ;
        RECT  -37.8 172.35 -36.9 173.25 ;
        RECT  -32.25 229.95 -7.95 230.85 ;
        RECT  -37.35 172.35 -7.95 173.25 ;
        RECT  -8.55 229.8 -7.35 231.0 ;
        RECT  -8.55 172.05 -7.35 173.25 ;
        RECT  -37.95 172.2 -36.75 173.4 ;
        RECT  -46.65 292.65 -45.45 293.85 ;
        RECT  -43.2 267.0 -42.3 267.9 ;
        RECT  -43.2 277.5 -42.3 278.4 ;
        RECT  -42.75 267.0 -36.9 267.9 ;
        RECT  -51.75 277.65 -42.75 278.55 ;
        RECT  -43.35 266.85 -42.15 268.05 ;
        RECT  -43.35 277.35 -42.15 278.55 ;
        RECT  -45.9 316.5 -45.0 317.4 ;
        RECT  -51.75 316.65 -45.45 317.55 ;
        RECT  -46.05 316.35 -44.85 317.55 ;
        RECT  -43.2 267.0 -42.3 267.9 ;
        RECT  -43.2 253.5 -42.3 254.4 ;
        RECT  -42.75 267.0 -36.9 267.9 ;
        RECT  -51.75 253.65 -42.75 254.55 ;
        RECT  -43.35 266.85 -42.15 268.05 ;
        RECT  -43.35 253.35 -42.15 254.55 ;
        RECT  -45.9 344.7 -45.0 345.6 ;
        RECT  -56.85 344.85 -45.45 345.75 ;
        RECT  -46.05 344.55 -44.85 345.75 ;
        RECT  -62.4 229.95 -61.5 230.85 ;
        RECT  -61.95 229.95 -22.65 230.85 ;
        RECT  -62.55 229.8 -61.35 231.0 ;
        RECT  -52.2 229.95 -51.3 230.85 ;
        RECT  -51.75 229.95 -22.65 230.85 ;
        RECT  -52.35 229.8 -51.15 231.0 ;
        RECT  -7.95 180.0 -7.05 189.6 ;
        RECT  -22.65 180.0 -21.75 189.6 ;
        RECT  -21.75 181.8 -19.35 183.0 ;
        RECT  -9.75 181.8 -7.95 183.0 ;
        RECT  -8.85 186.6 -7.95 187.8 ;
        RECT  -21.75 186.6 -20.55 187.8 ;
        RECT  -19.5 184.2 -10.05 185.4 ;
        RECT  -14.7 187.5 -13.8 189.6 ;
        RECT  -14.7 180.0 -13.8 184.2 ;
        RECT  -13.65 186.6 -12.45 187.8 ;
        RECT  -13.65 184.2 -12.45 185.4 ;
        RECT  -14.55 186.6 -13.35 187.8 ;
        RECT  -14.55 184.2 -13.35 185.4 ;
        RECT  -19.35 181.8 -18.15 183.0 ;
        RECT  -8.85 181.8 -7.65 183.0 ;
        RECT  -13.65 186.3 -12.45 187.5 ;
        RECT  -7.95 189.6 -7.05 199.2 ;
        RECT  -22.65 189.6 -21.75 199.2 ;
        RECT  -21.75 191.4 -19.35 192.6 ;
        RECT  -9.75 191.4 -7.95 192.6 ;
        RECT  -8.85 196.2 -7.95 197.4 ;
        RECT  -21.75 196.2 -20.55 197.4 ;
        RECT  -19.5 193.8 -10.05 195.0 ;
        RECT  -14.7 197.1 -13.8 199.2 ;
        RECT  -14.7 189.6 -13.8 193.8 ;
        RECT  -13.65 196.2 -12.45 197.4 ;
        RECT  -13.65 193.8 -12.45 195.0 ;
        RECT  -14.55 196.2 -13.35 197.4 ;
        RECT  -14.55 193.8 -13.35 195.0 ;
        RECT  -19.35 191.4 -18.15 192.6 ;
        RECT  -8.85 191.4 -7.65 192.6 ;
        RECT  -13.65 195.9 -12.45 197.1 ;
        RECT  -37.35 164.4 -36.45 180.0 ;
        RECT  -22.65 164.4 -21.75 180.0 ;
        RECT  -35.1 175.2 -24.0 176.1 ;
        RECT  -25.05 177.0 -22.2 177.9 ;
        RECT  -36.9 177.0 -33.3 177.9 ;
        RECT  -25.05 167.55 -22.2 168.45 ;
        RECT  -25.05 172.35 -22.2 173.25 ;
        RECT  -36.9 167.55 -34.05 168.45 ;
        RECT  -27.15 164.4 -26.25 168.6 ;
        RECT  -32.7 164.4 -31.8 166.5 ;
        RECT  -34.5 164.4 -33.6 166.5 ;
        RECT  -29.85 175.2 -28.95 180.0 ;
        RECT  -30.9 167.4 -28.2 168.6 ;
        RECT  -30.9 169.8 -28.2 171.0 ;
        RECT  -30.9 169.8 -28.2 171.0 ;
        RECT  -30.9 172.2 -28.2 173.4 ;
        RECT  -30.9 172.2 -28.2 173.4 ;
        RECT  -30.9 174.6 -28.2 175.8 ;
        RECT  -31.05 167.4 -29.85 168.6 ;
        RECT  -31.05 169.8 -29.85 171.0 ;
        RECT  -31.05 169.8 -29.85 171.0 ;
        RECT  -31.05 172.2 -29.85 173.4 ;
        RECT  -31.05 172.2 -29.85 173.4 ;
        RECT  -31.05 174.6 -29.85 175.8 ;
        RECT  -26.25 177.0 -25.05 178.2 ;
        RECT  -38.1 177.0 -35.4 178.2 ;
        RECT  -26.25 169.8 -25.05 171.0 ;
        RECT  -26.25 174.6 -25.05 175.8 ;
        RECT  -28.65 167.4 -27.45 168.6 ;
        RECT  -33.0 170.7 -31.8 171.9 ;
        RECT  -33.0 170.7 -31.8 171.9 ;
        RECT  -33.9 165.3 -32.7 166.5 ;
        RECT  -33.0 173.1 -31.8 174.3 ;
        RECT  -33.0 173.1 -31.8 174.3 ;
        RECT  -36.0 165.3 -34.8 166.5 ;
        RECT  -37.35 164.4 -36.45 180.0 ;
        RECT  -52.05 164.4 -51.15 180.0 ;
        RECT  -49.8 175.2 -38.7 176.1 ;
        RECT  -51.6 177.0 -48.75 177.9 ;
        RECT  -40.5 177.0 -36.9 177.9 ;
        RECT  -51.6 167.55 -48.75 168.45 ;
        RECT  -51.6 172.35 -48.75 173.25 ;
        RECT  -39.75 167.55 -36.9 168.45 ;
        RECT  -47.55 164.4 -46.65 168.6 ;
        RECT  -42.0 164.4 -41.1 166.5 ;
        RECT  -40.2 164.4 -39.3 166.5 ;
        RECT  -44.85 175.2 -43.95 180.0 ;
        RECT  -43.8 167.4 -41.1 168.6 ;
        RECT  -43.8 169.8 -41.1 171.0 ;
        RECT  -43.8 169.8 -41.1 171.0 ;
        RECT  -43.8 172.2 -41.1 173.4 ;
        RECT  -43.8 172.2 -41.1 173.4 ;
        RECT  -43.8 174.6 -41.1 175.8 ;
        RECT  -49.95 167.4 -48.75 168.6 ;
        RECT  -49.95 169.8 -48.75 171.0 ;
        RECT  -49.95 169.8 -48.75 171.0 ;
        RECT  -49.95 172.2 -48.75 173.4 ;
        RECT  -49.95 172.2 -48.75 173.4 ;
        RECT  -49.95 174.6 -48.75 175.8 ;
        RECT  -49.95 177.0 -48.75 178.2 ;
        RECT  -41.1 177.0 -38.4 178.2 ;
        RECT  -49.95 169.8 -48.75 171.0 ;
        RECT  -49.95 174.6 -48.75 175.8 ;
        RECT  -47.55 167.4 -46.35 168.6 ;
        RECT  -43.2 170.7 -42.0 171.9 ;
        RECT  -43.2 170.7 -42.0 171.9 ;
        RECT  -42.3 165.3 -41.1 166.5 ;
        RECT  -43.2 173.1 -42.0 174.3 ;
        RECT  -43.2 173.1 -42.0 174.3 ;
        RECT  -40.2 165.3 -39.0 166.5 ;
        RECT  -37.35 180.0 -36.45 189.6 ;
        RECT  -22.65 180.0 -21.75 189.6 ;
        RECT  -25.05 186.6 -22.65 187.8 ;
        RECT  -36.45 186.6 -34.65 187.8 ;
        RECT  -36.45 181.8 -35.55 183.0 ;
        RECT  -23.85 181.8 -22.65 183.0 ;
        RECT  -34.35 184.2 -24.9 185.4 ;
        RECT  -30.6 180.0 -29.7 182.1 ;
        RECT  -30.6 185.4 -29.7 189.6 ;
        RECT  -31.95 181.8 -30.75 183.0 ;
        RECT  -31.95 184.2 -30.75 185.4 ;
        RECT  -31.05 181.8 -29.85 183.0 ;
        RECT  -31.05 184.2 -29.85 185.4 ;
        RECT  -26.25 186.6 -25.05 187.8 ;
        RECT  -36.75 186.6 -35.55 187.8 ;
        RECT  -31.95 182.1 -30.75 183.3 ;
        RECT  -37.35 180.0 -36.45 189.6 ;
        RECT  -52.05 180.0 -51.15 189.6 ;
        RECT  -51.15 186.6 -48.75 187.8 ;
        RECT  -39.15 186.6 -37.35 187.8 ;
        RECT  -38.25 181.8 -37.35 183.0 ;
        RECT  -51.15 181.8 -49.95 183.0 ;
        RECT  -48.9 184.2 -39.45 185.4 ;
        RECT  -44.1 180.0 -43.2 182.1 ;
        RECT  -44.1 185.4 -43.2 189.6 ;
        RECT  -40.65 181.8 -39.45 183.0 ;
        RECT  -40.65 184.2 -39.45 185.4 ;
        RECT  -49.95 181.8 -48.75 183.0 ;
        RECT  -49.95 184.2 -48.75 185.4 ;
        RECT  -49.95 186.6 -48.75 187.8 ;
        RECT  -39.45 186.6 -38.25 187.8 ;
        RECT  -44.25 182.1 -43.05 183.3 ;
        RECT  -37.35 189.6 -36.45 199.2 ;
        RECT  -52.05 189.6 -51.15 199.2 ;
        RECT  -51.15 196.2 -48.75 197.4 ;
        RECT  -39.15 196.2 -37.35 197.4 ;
        RECT  -38.25 191.4 -37.35 192.6 ;
        RECT  -51.15 191.4 -49.95 192.6 ;
        RECT  -48.9 193.8 -39.45 195.0 ;
        RECT  -44.1 189.6 -43.2 191.7 ;
        RECT  -44.1 195.0 -43.2 199.2 ;
        RECT  -40.65 191.4 -39.45 192.6 ;
        RECT  -40.65 193.8 -39.45 195.0 ;
        RECT  -49.95 191.4 -48.75 192.6 ;
        RECT  -49.95 193.8 -48.75 195.0 ;
        RECT  -49.95 196.2 -48.75 197.4 ;
        RECT  -39.45 196.2 -38.25 197.4 ;
        RECT  -44.25 191.7 -43.05 192.9 ;
        RECT  -37.35 199.2 -36.45 208.8 ;
        RECT  -52.05 199.2 -51.15 208.8 ;
        RECT  -51.15 205.8 -48.75 207.0 ;
        RECT  -39.15 205.8 -37.35 207.0 ;
        RECT  -38.25 201.0 -37.35 202.2 ;
        RECT  -51.15 201.0 -49.95 202.2 ;
        RECT  -48.9 203.4 -39.45 204.6 ;
        RECT  -44.1 199.2 -43.2 201.3 ;
        RECT  -44.1 204.6 -43.2 208.8 ;
        RECT  -40.65 201.0 -39.45 202.2 ;
        RECT  -40.65 203.4 -39.45 204.6 ;
        RECT  -49.95 201.0 -48.75 202.2 ;
        RECT  -49.95 203.4 -48.75 204.6 ;
        RECT  -49.95 205.8 -48.75 207.0 ;
        RECT  -39.45 205.8 -38.25 207.0 ;
        RECT  -44.25 201.3 -43.05 202.5 ;
        RECT  -40.8 144.3 -39.6 145.5 ;
        RECT  -40.8 150.9 -39.6 152.1 ;
        RECT  -44.25 144.3 -43.05 145.5 ;
        RECT  -44.25 153.6 -43.05 154.8 ;
        RECT  -64.65 144.3 -63.45 145.5 ;
        RECT  -64.65 156.3 -63.45 157.5 ;
        RECT  -49.05 144.3 -47.85 145.5 ;
        RECT  -49.05 159.0 -47.85 160.2 ;
        RECT  -17.4 153.6 -16.2 154.8 ;
        RECT  -14.1 161.7 -12.9 162.9 ;
        RECT  -27.45 161.7 -26.25 162.9 ;
        RECT  -33.0 153.6 -31.8 154.8 ;
        RECT  -34.8 156.3 -33.6 157.5 ;
        RECT  -47.85 161.7 -46.65 162.9 ;
        RECT  -42.3 159.0 -41.1 160.2 ;
        RECT  -40.5 156.3 -39.3 157.5 ;
        RECT  -16.05 121.05 -15.15 121.95 ;
        RECT  -5.85 121.05 -4.95 121.95 ;
        RECT  -5.7 150.9 -4.8 151.8 ;
        RECT  -16.05 119.7 -15.15 121.5 ;
        RECT  -5.7 121.5 -4.8 151.35 ;
        RECT  -16.2 120.9 -15.0 122.1 ;
        RECT  -6.0 120.9 -4.8 122.1 ;
        RECT  -5.85 150.75 -4.65 151.95 ;
        RECT  -14.7 145.95 -13.8 146.85 ;
        RECT  -13.8 145.95 -12.9 146.85 ;
        RECT  -14.7 145.5 -13.8 146.4 ;
        RECT  -14.25 145.95 -13.35 146.85 ;
        RECT  -13.8 146.4 -12.9 164.4 ;
        RECT  -30.9 214.2 -29.7 215.4 ;
        RECT  -44.4 211.5 -43.2 212.7 ;
        RECT  -15.0 216.9 -13.8 218.1 ;
        RECT  -4.05 214.2 -3.15 215.1 ;
        RECT  -3.9 214.65 -3.0 265.2 ;
        RECT  -4.2 214.05 -3.0 215.25 ;
        RECT  -22.95 219.6 -21.75 220.8 ;
        RECT  -52.35 219.6 -51.15 220.8 ;
        RECT  -8.25 148.2 -7.05 149.4 ;
        RECT  -14.7 126.45 -13.8 127.35 ;
        RECT  -27.75 126.45 -26.85 127.35 ;
        RECT  -14.7 126.9 -13.8 128.7 ;
        RECT  -27.6 85.5 -26.7 126.9 ;
        RECT  -14.85 126.3 -13.65 127.5 ;
        RECT  -27.9 126.3 -26.7 127.5 ;
        RECT  -14.7 123.75 -13.8 124.65 ;
        RECT  -14.1 123.75 -13.2 124.65 ;
        RECT  -14.7 124.2 -13.8 126.9 ;
        RECT  -14.25 123.75 -13.65 124.65 ;
        RECT  -14.1 119.7 -13.2 124.2 ;
        RECT  -27.6 85.5 -26.4 86.7 ;
        RECT  -14.1 88.5 -12.9 89.7 ;
        RECT  -15.0 175.5 -13.8 176.7 ;
        RECT  -15.0 180.0 -13.8 181.2 ;
        RECT  0.0 219.6 2.4 220.8 ;
        Layer  via1 ; 
        RECT  124.8 209.7 125.4 210.3 ;
        RECT  133.8 209.7 134.4 210.3 ;
        RECT  125.7 200.4 126.3 201.0 ;
        RECT  129.9 200.4 130.5 201.0 ;
        RECT  124.8 219.3 125.4 219.9 ;
        RECT  133.8 219.3 134.4 219.9 ;
        RECT  125.7 228.6 126.3 229.2 ;
        RECT  129.9 228.6 130.5 229.2 ;
        RECT  124.8 239.1 125.4 239.7 ;
        RECT  133.8 239.1 134.4 239.7 ;
        RECT  125.7 229.8 126.3 230.4 ;
        RECT  129.9 229.8 130.5 230.4 ;
        RECT  124.8 248.7 125.4 249.3 ;
        RECT  133.8 248.7 134.4 249.3 ;
        RECT  125.7 258.0 126.3 258.6 ;
        RECT  129.9 258.0 130.5 258.6 ;
        RECT  124.8 268.5 125.4 269.1 ;
        RECT  133.8 268.5 134.4 269.1 ;
        RECT  125.7 259.2 126.3 259.8 ;
        RECT  129.9 259.2 130.5 259.8 ;
        RECT  124.8 278.1 125.4 278.7 ;
        RECT  133.8 278.1 134.4 278.7 ;
        RECT  125.7 287.4 126.3 288.0 ;
        RECT  129.9 287.4 130.5 288.0 ;
        RECT  124.8 297.9 125.4 298.5 ;
        RECT  133.8 297.9 134.4 298.5 ;
        RECT  125.7 288.6 126.3 289.2 ;
        RECT  129.9 288.6 130.5 289.2 ;
        RECT  124.8 307.5 125.4 308.1 ;
        RECT  133.8 307.5 134.4 308.1 ;
        RECT  125.7 316.8 126.3 317.4 ;
        RECT  129.9 316.8 130.5 317.4 ;
        RECT  124.8 327.3 125.4 327.9 ;
        RECT  133.8 327.3 134.4 327.9 ;
        RECT  125.7 318.0 126.3 318.6 ;
        RECT  129.9 318.0 130.5 318.6 ;
        RECT  124.8 336.9 125.4 337.5 ;
        RECT  133.8 336.9 134.4 337.5 ;
        RECT  125.7 346.2 126.3 346.8 ;
        RECT  129.9 346.2 130.5 346.8 ;
        RECT  124.8 356.7 125.4 357.3 ;
        RECT  133.8 356.7 134.4 357.3 ;
        RECT  125.7 347.4 126.3 348.0 ;
        RECT  129.9 347.4 130.5 348.0 ;
        RECT  124.8 366.3 125.4 366.9 ;
        RECT  133.8 366.3 134.4 366.9 ;
        RECT  125.7 375.6 126.3 376.2 ;
        RECT  129.9 375.6 130.5 376.2 ;
        RECT  124.8 386.1 125.4 386.7 ;
        RECT  133.8 386.1 134.4 386.7 ;
        RECT  125.7 376.8 126.3 377.4 ;
        RECT  129.9 376.8 130.5 377.4 ;
        RECT  124.8 395.7 125.4 396.3 ;
        RECT  133.8 395.7 134.4 396.3 ;
        RECT  125.7 405.0 126.3 405.6 ;
        RECT  129.9 405.0 130.5 405.6 ;
        RECT  124.8 415.5 125.4 416.1 ;
        RECT  133.8 415.5 134.4 416.1 ;
        RECT  125.7 406.2 126.3 406.8 ;
        RECT  129.9 406.2 130.5 406.8 ;
        RECT  124.8 425.1 125.4 425.7 ;
        RECT  133.8 425.1 134.4 425.7 ;
        RECT  125.7 434.4 126.3 435.0 ;
        RECT  129.9 434.4 130.5 435.0 ;
        RECT  135.0 209.7 135.6 210.3 ;
        RECT  144.0 209.7 144.6 210.3 ;
        RECT  135.9 200.4 136.5 201.0 ;
        RECT  140.1 200.4 140.7 201.0 ;
        RECT  135.0 219.3 135.6 219.9 ;
        RECT  144.0 219.3 144.6 219.9 ;
        RECT  135.9 228.6 136.5 229.2 ;
        RECT  140.1 228.6 140.7 229.2 ;
        RECT  135.0 239.1 135.6 239.7 ;
        RECT  144.0 239.1 144.6 239.7 ;
        RECT  135.9 229.8 136.5 230.4 ;
        RECT  140.1 229.8 140.7 230.4 ;
        RECT  135.0 248.7 135.6 249.3 ;
        RECT  144.0 248.7 144.6 249.3 ;
        RECT  135.9 258.0 136.5 258.6 ;
        RECT  140.1 258.0 140.7 258.6 ;
        RECT  135.0 268.5 135.6 269.1 ;
        RECT  144.0 268.5 144.6 269.1 ;
        RECT  135.9 259.2 136.5 259.8 ;
        RECT  140.1 259.2 140.7 259.8 ;
        RECT  135.0 278.1 135.6 278.7 ;
        RECT  144.0 278.1 144.6 278.7 ;
        RECT  135.9 287.4 136.5 288.0 ;
        RECT  140.1 287.4 140.7 288.0 ;
        RECT  135.0 297.9 135.6 298.5 ;
        RECT  144.0 297.9 144.6 298.5 ;
        RECT  135.9 288.6 136.5 289.2 ;
        RECT  140.1 288.6 140.7 289.2 ;
        RECT  135.0 307.5 135.6 308.1 ;
        RECT  144.0 307.5 144.6 308.1 ;
        RECT  135.9 316.8 136.5 317.4 ;
        RECT  140.1 316.8 140.7 317.4 ;
        RECT  135.0 327.3 135.6 327.9 ;
        RECT  144.0 327.3 144.6 327.9 ;
        RECT  135.9 318.0 136.5 318.6 ;
        RECT  140.1 318.0 140.7 318.6 ;
        RECT  135.0 336.9 135.6 337.5 ;
        RECT  144.0 336.9 144.6 337.5 ;
        RECT  135.9 346.2 136.5 346.8 ;
        RECT  140.1 346.2 140.7 346.8 ;
        RECT  135.0 356.7 135.6 357.3 ;
        RECT  144.0 356.7 144.6 357.3 ;
        RECT  135.9 347.4 136.5 348.0 ;
        RECT  140.1 347.4 140.7 348.0 ;
        RECT  135.0 366.3 135.6 366.9 ;
        RECT  144.0 366.3 144.6 366.9 ;
        RECT  135.9 375.6 136.5 376.2 ;
        RECT  140.1 375.6 140.7 376.2 ;
        RECT  135.0 386.1 135.6 386.7 ;
        RECT  144.0 386.1 144.6 386.7 ;
        RECT  135.9 376.8 136.5 377.4 ;
        RECT  140.1 376.8 140.7 377.4 ;
        RECT  135.0 395.7 135.6 396.3 ;
        RECT  144.0 395.7 144.6 396.3 ;
        RECT  135.9 405.0 136.5 405.6 ;
        RECT  140.1 405.0 140.7 405.6 ;
        RECT  135.0 415.5 135.6 416.1 ;
        RECT  144.0 415.5 144.6 416.1 ;
        RECT  135.9 406.2 136.5 406.8 ;
        RECT  140.1 406.2 140.7 406.8 ;
        RECT  135.0 425.1 135.6 425.7 ;
        RECT  144.0 425.1 144.6 425.7 ;
        RECT  135.9 434.4 136.5 435.0 ;
        RECT  140.1 434.4 140.7 435.0 ;
        RECT  145.2 209.7 145.8 210.3 ;
        RECT  154.2 209.7 154.8 210.3 ;
        RECT  146.1 200.4 146.7 201.0 ;
        RECT  150.3 200.4 150.9 201.0 ;
        RECT  145.2 219.3 145.8 219.9 ;
        RECT  154.2 219.3 154.8 219.9 ;
        RECT  146.1 228.6 146.7 229.2 ;
        RECT  150.3 228.6 150.9 229.2 ;
        RECT  145.2 239.1 145.8 239.7 ;
        RECT  154.2 239.1 154.8 239.7 ;
        RECT  146.1 229.8 146.7 230.4 ;
        RECT  150.3 229.8 150.9 230.4 ;
        RECT  145.2 248.7 145.8 249.3 ;
        RECT  154.2 248.7 154.8 249.3 ;
        RECT  146.1 258.0 146.7 258.6 ;
        RECT  150.3 258.0 150.9 258.6 ;
        RECT  145.2 268.5 145.8 269.1 ;
        RECT  154.2 268.5 154.8 269.1 ;
        RECT  146.1 259.2 146.7 259.8 ;
        RECT  150.3 259.2 150.9 259.8 ;
        RECT  145.2 278.1 145.8 278.7 ;
        RECT  154.2 278.1 154.8 278.7 ;
        RECT  146.1 287.4 146.7 288.0 ;
        RECT  150.3 287.4 150.9 288.0 ;
        RECT  145.2 297.9 145.8 298.5 ;
        RECT  154.2 297.9 154.8 298.5 ;
        RECT  146.1 288.6 146.7 289.2 ;
        RECT  150.3 288.6 150.9 289.2 ;
        RECT  145.2 307.5 145.8 308.1 ;
        RECT  154.2 307.5 154.8 308.1 ;
        RECT  146.1 316.8 146.7 317.4 ;
        RECT  150.3 316.8 150.9 317.4 ;
        RECT  145.2 327.3 145.8 327.9 ;
        RECT  154.2 327.3 154.8 327.9 ;
        RECT  146.1 318.0 146.7 318.6 ;
        RECT  150.3 318.0 150.9 318.6 ;
        RECT  145.2 336.9 145.8 337.5 ;
        RECT  154.2 336.9 154.8 337.5 ;
        RECT  146.1 346.2 146.7 346.8 ;
        RECT  150.3 346.2 150.9 346.8 ;
        RECT  145.2 356.7 145.8 357.3 ;
        RECT  154.2 356.7 154.8 357.3 ;
        RECT  146.1 347.4 146.7 348.0 ;
        RECT  150.3 347.4 150.9 348.0 ;
        RECT  145.2 366.3 145.8 366.9 ;
        RECT  154.2 366.3 154.8 366.9 ;
        RECT  146.1 375.6 146.7 376.2 ;
        RECT  150.3 375.6 150.9 376.2 ;
        RECT  145.2 386.1 145.8 386.7 ;
        RECT  154.2 386.1 154.8 386.7 ;
        RECT  146.1 376.8 146.7 377.4 ;
        RECT  150.3 376.8 150.9 377.4 ;
        RECT  145.2 395.7 145.8 396.3 ;
        RECT  154.2 395.7 154.8 396.3 ;
        RECT  146.1 405.0 146.7 405.6 ;
        RECT  150.3 405.0 150.9 405.6 ;
        RECT  145.2 415.5 145.8 416.1 ;
        RECT  154.2 415.5 154.8 416.1 ;
        RECT  146.1 406.2 146.7 406.8 ;
        RECT  150.3 406.2 150.9 406.8 ;
        RECT  145.2 425.1 145.8 425.7 ;
        RECT  154.2 425.1 154.8 425.7 ;
        RECT  146.1 434.4 146.7 435.0 ;
        RECT  150.3 434.4 150.9 435.0 ;
        RECT  127.2 451.2 127.8 451.8 ;
        RECT  132.0 451.2 132.6 451.8 ;
        RECT  127.2 442.8 127.8 443.4 ;
        RECT  129.6 442.8 130.2 443.4 ;
        RECT  137.4 451.2 138.0 451.8 ;
        RECT  142.2 451.2 142.8 451.8 ;
        RECT  137.4 442.8 138.0 443.4 ;
        RECT  139.8 442.8 140.4 443.4 ;
        RECT  147.6 451.2 148.2 451.8 ;
        RECT  152.4 451.2 153.0 451.8 ;
        RECT  147.6 442.8 148.2 443.4 ;
        RECT  150.0 442.8 150.6 443.4 ;
        RECT  133.8 194.1 134.4 194.7 ;
        RECT  128.1 164.7 128.7 165.3 ;
        RECT  130.8 164.7 131.4 165.3 ;
        RECT  125.1 154.8 125.7 155.4 ;
        RECT  144.0 194.1 144.6 194.7 ;
        RECT  138.3 164.7 138.9 165.3 ;
        RECT  141.0 164.7 141.6 165.3 ;
        RECT  135.3 154.8 135.9 155.4 ;
        RECT  154.2 194.1 154.8 194.7 ;
        RECT  148.5 164.7 149.1 165.3 ;
        RECT  151.2 164.7 151.8 165.3 ;
        RECT  145.5 154.8 146.1 155.4 ;
        RECT  125.7 148.2 126.3 148.8 ;
        RECT  130.2 147.6 130.8 148.2 ;
        RECT  127.5 138.0 128.1 138.6 ;
        RECT  126.6 126.3 127.2 126.9 ;
        RECT  133.2 115.5 133.8 116.1 ;
        RECT  129.9 110.1 130.5 110.7 ;
        RECT  126.6 100.2 127.2 100.8 ;
        RECT  133.8 96.0 134.4 96.6 ;
        RECT  127.8 93.9 128.4 94.5 ;
        RECT  135.9 148.2 136.5 148.8 ;
        RECT  140.4 147.6 141.0 148.2 ;
        RECT  137.7 138.0 138.3 138.6 ;
        RECT  136.8 126.3 137.4 126.9 ;
        RECT  143.4 115.5 144.0 116.1 ;
        RECT  140.1 110.1 140.7 110.7 ;
        RECT  136.8 100.2 137.4 100.8 ;
        RECT  144.0 96.0 144.6 96.6 ;
        RECT  138.0 93.9 138.6 94.5 ;
        RECT  146.1 148.2 146.7 148.8 ;
        RECT  150.6 147.6 151.2 148.2 ;
        RECT  147.9 138.0 148.5 138.6 ;
        RECT  147.0 126.3 147.6 126.9 ;
        RECT  153.6 115.5 154.2 116.1 ;
        RECT  150.3 110.1 150.9 110.7 ;
        RECT  147.0 100.2 147.6 100.8 ;
        RECT  154.2 96.0 154.8 96.6 ;
        RECT  148.2 93.9 148.8 94.5 ;
        RECT  127.8 85.5 128.4 86.1 ;
        RECT  130.2 81.0 130.8 81.6 ;
        RECT  129.3 77.7 129.9 78.3 ;
        RECT  133.8 77.1 134.4 77.7 ;
        RECT  129.3 75.6 129.9 76.2 ;
        RECT  126.0 74.7 126.6 75.3 ;
        RECT  130.2 71.1 130.8 71.7 ;
        RECT  130.2 68.7 130.8 69.3 ;
        RECT  127.8 65.7 128.4 66.3 ;
        RECT  128.7 62.4 129.3 63.0 ;
        RECT  126.0 61.2 126.6 61.8 ;
        RECT  130.2 55.5 130.8 56.1 ;
        RECT  129.3 52.2 129.9 52.8 ;
        RECT  133.8 51.6 134.4 52.2 ;
        RECT  129.3 49.2 129.9 49.8 ;
        RECT  126.0 48.3 126.6 48.9 ;
        RECT  130.2 44.7 130.8 45.3 ;
        RECT  130.2 42.3 130.8 42.9 ;
        RECT  127.8 39.3 128.4 39.9 ;
        RECT  139.8 85.5 140.4 86.1 ;
        RECT  137.4 81.0 138.0 81.6 ;
        RECT  138.3 77.7 138.9 78.3 ;
        RECT  133.8 77.1 134.4 77.7 ;
        RECT  138.3 75.6 138.9 76.2 ;
        RECT  141.6 74.7 142.2 75.3 ;
        RECT  137.4 71.1 138.0 71.7 ;
        RECT  137.4 68.7 138.0 69.3 ;
        RECT  139.8 65.7 140.4 66.3 ;
        RECT  138.9 62.4 139.5 63.0 ;
        RECT  141.6 61.2 142.2 61.8 ;
        RECT  137.4 55.5 138.0 56.1 ;
        RECT  138.3 52.2 138.9 52.8 ;
        RECT  133.8 51.6 134.4 52.2 ;
        RECT  138.3 49.2 138.9 49.8 ;
        RECT  141.6 48.3 142.2 48.9 ;
        RECT  137.4 44.7 138.0 45.3 ;
        RECT  137.4 42.3 138.0 42.9 ;
        RECT  139.8 39.3 140.4 39.9 ;
        RECT  148.2 85.5 148.8 86.1 ;
        RECT  150.6 81.0 151.2 81.6 ;
        RECT  149.7 77.7 150.3 78.3 ;
        RECT  154.2 77.1 154.8 77.7 ;
        RECT  149.7 75.6 150.3 76.2 ;
        RECT  146.4 74.7 147.0 75.3 ;
        RECT  150.6 71.1 151.2 71.7 ;
        RECT  150.6 68.7 151.2 69.3 ;
        RECT  148.2 65.7 148.8 66.3 ;
        RECT  149.1 62.4 149.7 63.0 ;
        RECT  146.4 61.2 147.0 61.8 ;
        RECT  150.6 55.5 151.2 56.1 ;
        RECT  149.7 52.2 150.3 52.8 ;
        RECT  154.2 51.6 154.8 52.2 ;
        RECT  149.7 49.2 150.3 49.8 ;
        RECT  146.4 48.3 147.0 48.9 ;
        RECT  150.6 44.7 151.2 45.3 ;
        RECT  150.6 42.3 151.2 42.9 ;
        RECT  148.2 39.3 148.8 39.9 ;
        RECT  126.9 45.0 127.5 45.6 ;
        RECT  131.7 41.4 132.3 42.0 ;
        RECT  133.8 36.9 134.4 37.5 ;
        RECT  140.7 45.0 141.3 45.6 ;
        RECT  135.9 41.4 136.5 42.0 ;
        RECT  133.8 36.9 134.4 37.5 ;
        RECT  147.3 45.0 147.9 45.6 ;
        RECT  152.1 41.4 152.7 42.0 ;
        RECT  154.2 36.9 154.8 37.5 ;
        RECT  58.5 93.15 59.1 93.75 ;
        RECT  77.7 87.9 78.3 88.5 ;
        RECT  56.4 98.55 57.0 99.15 ;
        RECT  75.6 103.8 76.2 104.4 ;
        RECT  58.5 90.3 59.1 90.9 ;
        RECT  56.4 87.0 57.0 87.6 ;
        RECT  54.3 101.4 54.9 102.0 ;
        RECT  56.4 104.7 57.0 105.3 ;
        RECT  58.5 119.7 59.1 120.3 ;
        RECT  52.2 116.4 52.8 117.0 ;
        RECT  54.3 130.8 54.9 131.4 ;
        RECT  77.7 130.8 78.3 131.4 ;
        RECT  52.2 134.1 52.8 134.7 ;
        RECT  75.6 134.1 76.2 134.7 ;
        RECT  60.6 81.15 61.2 81.75 ;
        RECT  62.7 95.85 63.3 96.45 ;
        RECT  60.6 110.55 61.2 111.15 ;
        RECT  62.7 125.25 63.3 125.85 ;
        RECT  60.6 137.7 61.2 138.3 ;
        RECT  58.5 151.95 59.1 152.55 ;
        RECT  77.7 146.7 78.3 147.3 ;
        RECT  56.4 157.35 57.0 157.95 ;
        RECT  75.6 162.6 76.2 163.2 ;
        RECT  58.5 149.1 59.1 149.7 ;
        RECT  56.4 145.8 57.0 146.4 ;
        RECT  54.3 160.2 54.9 160.8 ;
        RECT  56.4 163.5 57.0 164.1 ;
        RECT  58.5 178.5 59.1 179.1 ;
        RECT  52.2 175.2 52.8 175.8 ;
        RECT  54.3 189.6 54.9 190.2 ;
        RECT  77.7 189.6 78.3 190.2 ;
        RECT  52.2 192.9 52.8 193.5 ;
        RECT  75.6 192.9 76.2 193.5 ;
        RECT  60.6 139.95 61.2 140.55 ;
        RECT  62.7 154.65 63.3 155.25 ;
        RECT  60.6 169.35 61.2 169.95 ;
        RECT  62.7 184.05 63.3 184.65 ;
        RECT  60.6 196.5 61.2 197.1 ;
        RECT  12.9 89.1 13.5 89.7 ;
        RECT  15.0 105.0 15.6 105.6 ;
        RECT  17.1 118.5 17.7 119.1 ;
        RECT  19.2 134.4 19.8 135.0 ;
        RECT  21.3 147.9 21.9 148.5 ;
        RECT  23.4 163.8 24.0 164.4 ;
        RECT  25.5 177.3 26.1 177.9 ;
        RECT  27.6 193.2 28.2 193.8 ;
        RECT  12.9 209.1 13.5 209.7 ;
        RECT  21.3 205.8 21.9 206.4 ;
        RECT  12.9 220.2 13.5 220.8 ;
        RECT  23.4 223.5 24.0 224.1 ;
        RECT  12.9 238.5 13.5 239.1 ;
        RECT  25.5 235.2 26.1 235.8 ;
        RECT  12.9 249.6 13.5 250.2 ;
        RECT  27.6 252.9 28.2 253.5 ;
        RECT  15.0 267.9 15.6 268.5 ;
        RECT  21.3 264.6 21.9 265.2 ;
        RECT  15.0 279.0 15.6 279.6 ;
        RECT  23.4 282.3 24.0 282.9 ;
        RECT  15.0 297.3 15.6 297.9 ;
        RECT  25.5 294.0 26.1 294.6 ;
        RECT  15.0 308.4 15.6 309.0 ;
        RECT  27.6 311.7 28.2 312.3 ;
        RECT  17.1 326.7 17.7 327.3 ;
        RECT  21.3 323.4 21.9 324.0 ;
        RECT  17.1 337.8 17.7 338.4 ;
        RECT  23.4 341.1 24.0 341.7 ;
        RECT  17.1 356.1 17.7 356.7 ;
        RECT  25.5 352.8 26.1 353.4 ;
        RECT  17.1 367.2 17.7 367.8 ;
        RECT  27.6 370.5 28.2 371.1 ;
        RECT  19.2 385.5 19.8 386.1 ;
        RECT  21.3 382.2 21.9 382.8 ;
        RECT  19.2 396.6 19.8 397.2 ;
        RECT  23.4 399.9 24.0 400.5 ;
        RECT  19.2 414.9 19.8 415.5 ;
        RECT  25.5 411.6 26.1 412.2 ;
        RECT  19.2 426.0 19.8 426.6 ;
        RECT  27.6 429.3 28.2 429.9 ;
        RECT  51.0 214.65 51.6 215.25 ;
        RECT  57.3 214.65 57.9 215.25 ;
        RECT  67.2 209.1 67.8 209.7 ;
        RECT  51.3 209.1 51.9 209.7 ;
        RECT  51.0 229.35 51.6 229.95 ;
        RECT  57.3 229.35 57.9 229.95 ;
        RECT  67.2 219.9 67.8 220.5 ;
        RECT  51.3 219.9 51.9 220.5 ;
        RECT  51.0 244.05 51.6 244.65 ;
        RECT  57.3 244.05 57.9 244.65 ;
        RECT  67.2 238.5 67.8 239.1 ;
        RECT  51.3 238.5 51.9 239.1 ;
        RECT  51.0 258.75 51.6 259.35 ;
        RECT  57.3 258.75 57.9 259.35 ;
        RECT  67.2 249.3 67.8 249.9 ;
        RECT  51.3 249.3 51.9 249.9 ;
        RECT  51.0 273.45 51.6 274.05 ;
        RECT  57.3 273.45 57.9 274.05 ;
        RECT  67.2 267.9 67.8 268.5 ;
        RECT  51.3 267.9 51.9 268.5 ;
        RECT  51.0 288.15 51.6 288.75 ;
        RECT  57.3 288.15 57.9 288.75 ;
        RECT  67.2 278.7 67.8 279.3 ;
        RECT  51.3 278.7 51.9 279.3 ;
        RECT  51.0 302.85 51.6 303.45 ;
        RECT  57.3 302.85 57.9 303.45 ;
        RECT  67.2 297.3 67.8 297.9 ;
        RECT  51.3 297.3 51.9 297.9 ;
        RECT  51.0 317.55 51.6 318.15 ;
        RECT  57.3 317.55 57.9 318.15 ;
        RECT  67.2 308.1 67.8 308.7 ;
        RECT  51.3 308.1 51.9 308.7 ;
        RECT  51.0 332.25 51.6 332.85 ;
        RECT  57.3 332.25 57.9 332.85 ;
        RECT  67.2 326.7 67.8 327.3 ;
        RECT  51.3 326.7 51.9 327.3 ;
        RECT  51.0 346.95 51.6 347.55 ;
        RECT  57.3 346.95 57.9 347.55 ;
        RECT  67.2 337.5 67.8 338.1 ;
        RECT  51.3 337.5 51.9 338.1 ;
        RECT  51.0 361.65 51.6 362.25 ;
        RECT  57.3 361.65 57.9 362.25 ;
        RECT  67.2 356.1 67.8 356.7 ;
        RECT  51.3 356.1 51.9 356.7 ;
        RECT  51.0 376.35 51.6 376.95 ;
        RECT  57.3 376.35 57.9 376.95 ;
        RECT  67.2 366.9 67.8 367.5 ;
        RECT  51.3 366.9 51.9 367.5 ;
        RECT  51.0 391.05 51.6 391.65 ;
        RECT  57.3 391.05 57.9 391.65 ;
        RECT  67.2 385.5 67.8 386.1 ;
        RECT  51.3 385.5 51.9 386.1 ;
        RECT  51.0 405.75 51.6 406.35 ;
        RECT  57.3 405.75 57.9 406.35 ;
        RECT  67.2 396.3 67.8 396.9 ;
        RECT  51.3 396.3 51.9 396.9 ;
        RECT  51.0 420.45 51.6 421.05 ;
        RECT  57.3 420.45 57.9 421.05 ;
        RECT  67.2 414.9 67.8 415.5 ;
        RECT  51.3 414.9 51.9 415.5 ;
        RECT  51.0 435.15 51.6 435.75 ;
        RECT  57.3 435.15 57.9 435.75 ;
        RECT  67.2 425.7 67.8 426.3 ;
        RECT  51.3 425.7 51.9 426.3 ;
        RECT  69.9 75.3 70.5 75.9 ;
        RECT  65.4 72.9 66.0 73.5 ;
        RECT  62.1 73.8 62.7 74.4 ;
        RECT  61.5 69.3 62.1 69.9 ;
        RECT  60.0 73.8 60.6 74.4 ;
        RECT  59.1 77.1 59.7 77.7 ;
        RECT  55.5 72.9 56.1 73.5 ;
        RECT  53.1 72.9 53.7 73.5 ;
        RECT  50.1 75.3 50.7 75.9 ;
        RECT  46.8 74.4 47.4 75.0 ;
        RECT  45.6 77.1 46.2 77.7 ;
        RECT  39.9 72.9 40.5 73.5 ;
        RECT  36.6 73.8 37.2 74.4 ;
        RECT  36.0 69.3 36.6 69.9 ;
        RECT  33.6 73.8 34.2 74.4 ;
        RECT  32.7 77.1 33.3 77.7 ;
        RECT  29.1 72.9 29.7 73.5 ;
        RECT  26.7 72.9 27.3 73.5 ;
        RECT  23.7 75.3 24.3 75.9 ;
        RECT  69.9 63.3 70.5 63.9 ;
        RECT  65.4 65.7 66.0 66.3 ;
        RECT  62.1 64.8 62.7 65.4 ;
        RECT  61.5 69.3 62.1 69.9 ;
        RECT  60.0 64.8 60.6 65.4 ;
        RECT  59.1 61.5 59.7 62.1 ;
        RECT  55.5 65.7 56.1 66.3 ;
        RECT  53.1 65.7 53.7 66.3 ;
        RECT  50.1 63.3 50.7 63.9 ;
        RECT  46.8 64.2 47.4 64.8 ;
        RECT  45.6 61.5 46.2 62.1 ;
        RECT  39.9 65.7 40.5 66.3 ;
        RECT  36.6 64.8 37.2 65.4 ;
        RECT  36.0 69.3 36.6 69.9 ;
        RECT  33.6 64.8 34.2 65.4 ;
        RECT  32.7 61.5 33.3 62.1 ;
        RECT  29.1 65.7 29.7 66.3 ;
        RECT  26.7 65.7 27.3 66.3 ;
        RECT  23.7 63.3 24.3 63.9 ;
        RECT  69.9 54.9 70.5 55.5 ;
        RECT  65.4 52.5 66.0 53.1 ;
        RECT  62.1 53.4 62.7 54.0 ;
        RECT  61.5 48.9 62.1 49.5 ;
        RECT  60.0 53.4 60.6 54.0 ;
        RECT  59.1 56.7 59.7 57.3 ;
        RECT  55.5 52.5 56.1 53.1 ;
        RECT  53.1 52.5 53.7 53.1 ;
        RECT  50.1 54.9 50.7 55.5 ;
        RECT  46.8 54.0 47.4 54.6 ;
        RECT  45.6 56.7 46.2 57.3 ;
        RECT  39.9 52.5 40.5 53.1 ;
        RECT  36.6 53.4 37.2 54.0 ;
        RECT  36.0 48.9 36.6 49.5 ;
        RECT  33.6 53.4 34.2 54.0 ;
        RECT  32.7 56.7 33.3 57.3 ;
        RECT  29.1 52.5 29.7 53.1 ;
        RECT  26.7 52.5 27.3 53.1 ;
        RECT  23.7 54.9 24.3 55.5 ;
        RECT  69.9 42.9 70.5 43.5 ;
        RECT  65.4 45.3 66.0 45.9 ;
        RECT  62.1 44.4 62.7 45.0 ;
        RECT  61.5 48.9 62.1 49.5 ;
        RECT  60.0 44.4 60.6 45.0 ;
        RECT  59.1 41.1 59.7 41.7 ;
        RECT  55.5 45.3 56.1 45.9 ;
        RECT  53.1 45.3 53.7 45.9 ;
        RECT  50.1 42.9 50.7 43.5 ;
        RECT  46.8 43.8 47.4 44.4 ;
        RECT  45.6 41.1 46.2 41.7 ;
        RECT  39.9 45.3 40.5 45.9 ;
        RECT  36.6 44.4 37.2 45.0 ;
        RECT  36.0 48.9 36.6 49.5 ;
        RECT  33.6 44.4 34.2 45.0 ;
        RECT  32.7 41.1 33.3 41.7 ;
        RECT  29.1 45.3 29.7 45.9 ;
        RECT  26.7 45.3 27.3 45.9 ;
        RECT  23.7 42.9 24.3 43.5 ;
        RECT  90.9 89.1 91.5 89.7 ;
        RECT  88.2 105.0 88.8 105.6 ;
        RECT  85.5 147.9 86.1 148.5 ;
        RECT  82.8 163.8 83.4 164.4 ;
        RECT  114.3 33.6 114.9 34.2 ;
        RECT  108.9 28.95 109.5 29.55 ;
        RECT  111.6 26.55 112.2 27.15 ;
        RECT  114.3 446.7 114.9 447.3 ;
        RECT  117.0 98.25 117.6 98.85 ;
        RECT  119.7 196.35 120.3 196.95 ;
        RECT  16.8 76.8 17.4 77.4 ;
        RECT  106.2 456.9 106.8 457.5 ;
        RECT  95.4 437.4 96.0 438.0 ;
        RECT  96.6 437.4 97.2 438.0 ;
        RECT  134.1 437.4 134.7 438.0 ;
        RECT  144.3 437.4 144.9 438.0 ;
        RECT  154.5 437.4 155.1 438.0 ;
        RECT  123.0 437.4 123.6 438.0 ;
        RECT  102.0 8.4 102.6 9.0 ;
        RECT  103.2 8.4 103.8 9.0 ;
        RECT  133.8 8.4 134.4 9.0 ;
        RECT  133.8 8.4 134.4 9.0 ;
        RECT  154.2 8.4 154.8 9.0 ;
        RECT  88.05 229.35 88.65 229.95 ;
        RECT  88.05 258.75 88.65 259.35 ;
        RECT  88.05 288.15 88.65 288.75 ;
        RECT  88.05 317.55 88.65 318.15 ;
        RECT  88.05 346.95 88.65 347.55 ;
        RECT  88.05 376.35 88.65 376.95 ;
        RECT  88.05 405.75 88.65 406.35 ;
        RECT  88.05 435.15 88.65 435.75 ;
        RECT  95.4 140.85 96.0 141.45 ;
        RECT  96.6 140.85 97.2 141.45 ;
        RECT  95.4 199.65 96.0 200.25 ;
        RECT  96.6 199.65 97.2 200.25 ;
        RECT  75.3 69.45 75.9 70.05 ;
        RECT  95.4 69.45 96.0 70.05 ;
        RECT  96.6 69.45 97.2 70.05 ;
        RECT  75.3 69.45 75.9 70.05 ;
        RECT  95.4 69.45 96.0 70.05 ;
        RECT  96.6 69.45 97.2 70.05 ;
        RECT  75.3 49.05 75.9 49.65 ;
        RECT  95.4 49.05 96.0 49.65 ;
        RECT  96.6 49.05 97.2 49.65 ;
        RECT  75.3 49.05 75.9 49.65 ;
        RECT  95.4 49.05 96.0 49.65 ;
        RECT  96.6 49.05 97.2 49.65 ;
        RECT  -62.4 140.1 -61.8 140.7 ;
        RECT  -60.0 135.6 -59.4 136.2 ;
        RECT  -60.9 132.3 -60.3 132.9 ;
        RECT  -56.4 131.7 -55.8 132.3 ;
        RECT  -60.9 130.2 -60.3 130.8 ;
        RECT  -64.2 129.3 -63.6 129.9 ;
        RECT  -60.0 125.7 -59.4 126.3 ;
        RECT  -60.0 123.3 -59.4 123.9 ;
        RECT  -62.4 120.3 -61.8 120.9 ;
        RECT  -61.5 117.0 -60.9 117.6 ;
        RECT  -64.2 115.8 -63.6 116.4 ;
        RECT  -60.0 110.1 -59.4 110.7 ;
        RECT  -60.9 106.8 -60.3 107.4 ;
        RECT  -56.4 106.2 -55.8 106.8 ;
        RECT  -60.9 103.8 -60.3 104.4 ;
        RECT  -64.2 102.9 -63.6 103.5 ;
        RECT  -60.0 99.3 -59.4 99.9 ;
        RECT  -60.0 96.9 -59.4 97.5 ;
        RECT  -62.4 93.9 -61.8 94.5 ;
        RECT  -50.4 140.1 -49.8 140.7 ;
        RECT  -52.8 135.6 -52.2 136.2 ;
        RECT  -51.9 132.3 -51.3 132.9 ;
        RECT  -56.4 131.7 -55.8 132.3 ;
        RECT  -51.9 130.2 -51.3 130.8 ;
        RECT  -48.6 129.3 -48.0 129.9 ;
        RECT  -52.8 125.7 -52.2 126.3 ;
        RECT  -52.8 123.3 -52.2 123.9 ;
        RECT  -50.4 120.3 -49.8 120.9 ;
        RECT  -51.3 117.0 -50.7 117.6 ;
        RECT  -48.6 115.8 -48.0 116.4 ;
        RECT  -52.8 110.1 -52.2 110.7 ;
        RECT  -51.9 106.8 -51.3 107.4 ;
        RECT  -56.4 106.2 -55.8 106.8 ;
        RECT  -51.9 103.8 -51.3 104.4 ;
        RECT  -48.6 102.9 -48.0 103.5 ;
        RECT  -52.8 99.3 -52.2 99.9 ;
        RECT  -52.8 96.9 -52.2 97.5 ;
        RECT  -50.4 93.9 -49.8 94.5 ;
        RECT  -42.0 140.1 -41.4 140.7 ;
        RECT  -39.6 135.6 -39.0 136.2 ;
        RECT  -40.5 132.3 -39.9 132.9 ;
        RECT  -36.0 131.7 -35.4 132.3 ;
        RECT  -40.5 130.2 -39.9 130.8 ;
        RECT  -43.8 129.3 -43.2 129.9 ;
        RECT  -39.6 125.7 -39.0 126.3 ;
        RECT  -39.6 123.3 -39.0 123.9 ;
        RECT  -42.0 120.3 -41.4 120.9 ;
        RECT  -41.1 117.0 -40.5 117.6 ;
        RECT  -43.8 115.8 -43.2 116.4 ;
        RECT  -39.6 110.1 -39.0 110.7 ;
        RECT  -40.5 106.8 -39.9 107.4 ;
        RECT  -36.0 106.2 -35.4 106.8 ;
        RECT  -40.5 103.8 -39.9 104.4 ;
        RECT  -43.8 102.9 -43.2 103.5 ;
        RECT  -39.6 99.3 -39.0 99.9 ;
        RECT  -39.6 96.9 -39.0 97.5 ;
        RECT  -42.0 93.9 -41.4 94.5 ;
        RECT  -19.35 100.2 -18.75 100.8 ;
        RECT  -13.95 100.2 -13.35 100.8 ;
        RECT  -19.35 95.4 -18.75 96.0 ;
        RECT  -13.95 95.4 -13.35 96.0 ;
        RECT  -14.55 266.1 -13.95 266.7 ;
        RECT  -14.55 256.5 -13.95 257.1 ;
        RECT  -31.35 248.1 -30.75 248.7 ;
        RECT  -31.35 257.7 -30.75 258.3 ;
        RECT  -14.55 260.7 -13.95 261.3 ;
        RECT  -14.55 251.1 -13.95 251.7 ;
        RECT  -31.35 253.5 -30.75 254.1 ;
        RECT  -53.25 263.7 -52.65 264.3 ;
        RECT  -62.25 263.7 -61.65 264.3 ;
        RECT  -54.15 254.4 -53.55 255.0 ;
        RECT  -58.35 254.4 -57.75 255.0 ;
        RECT  -53.25 243.9 -52.65 244.5 ;
        RECT  -62.25 243.9 -61.65 244.5 ;
        RECT  -54.15 253.2 -53.55 253.8 ;
        RECT  -58.35 253.2 -57.75 253.8 ;
        RECT  -53.25 234.3 -52.65 234.9 ;
        RECT  -62.25 234.3 -61.65 234.9 ;
        RECT  -54.15 225.0 -53.55 225.6 ;
        RECT  -58.35 225.0 -57.75 225.6 ;
        RECT  -42.75 235.65 -42.15 236.25 ;
        RECT  -32.55 238.2 -31.95 238.8 ;
        RECT  -44.85 238.35 -44.25 238.95 ;
        RECT  -55.65 271.2 -55.05 271.8 ;
        RECT  -13.5 220.65 -12.9 221.25 ;
        RECT  -31.95 220.8 -31.35 221.4 ;
        RECT  -32.55 271.5 -31.95 272.1 ;
        RECT  -13.5 239.85 -12.9 240.45 ;
        RECT  -49.95 249.9 -49.35 250.5 ;
        RECT  -45.75 244.8 -45.15 245.4 ;
        RECT  -45.75 264.9 -45.15 265.5 ;
        RECT  -8.25 230.1 -7.65 230.7 ;
        RECT  -8.25 172.35 -7.65 172.95 ;
        RECT  -37.65 172.5 -37.05 173.1 ;
        RECT  -46.35 292.95 -45.75 293.55 ;
        RECT  -43.05 267.15 -42.45 267.75 ;
        RECT  -43.05 277.65 -42.45 278.25 ;
        RECT  -45.75 316.65 -45.15 317.25 ;
        RECT  -43.05 267.15 -42.45 267.75 ;
        RECT  -43.05 253.65 -42.45 254.25 ;
        RECT  -45.75 344.85 -45.15 345.45 ;
        RECT  -62.25 230.1 -61.65 230.7 ;
        RECT  -52.05 230.1 -51.45 230.7 ;
        RECT  -25.95 170.1 -25.35 170.7 ;
        RECT  -25.95 174.9 -25.35 175.5 ;
        RECT  -32.7 171.0 -32.1 171.6 ;
        RECT  -33.6 165.6 -33.0 166.2 ;
        RECT  -32.7 173.4 -32.1 174.0 ;
        RECT  -35.7 165.6 -35.1 166.2 ;
        RECT  -49.65 170.1 -49.05 170.7 ;
        RECT  -49.65 174.9 -49.05 175.5 ;
        RECT  -42.9 171.0 -42.3 171.6 ;
        RECT  -42.0 165.6 -41.4 166.2 ;
        RECT  -42.9 173.4 -42.3 174.0 ;
        RECT  -39.9 165.6 -39.3 166.2 ;
        RECT  -40.5 144.6 -39.9 145.2 ;
        RECT  -40.5 151.2 -39.9 151.8 ;
        RECT  -43.95 144.6 -43.35 145.2 ;
        RECT  -43.95 153.9 -43.35 154.5 ;
        RECT  -64.35 144.6 -63.75 145.2 ;
        RECT  -64.35 156.6 -63.75 157.2 ;
        RECT  -48.75 144.6 -48.15 145.2 ;
        RECT  -48.75 159.3 -48.15 159.9 ;
        RECT  -17.1 153.9 -16.5 154.5 ;
        RECT  -13.8 162.0 -13.2 162.6 ;
        RECT  -27.15 162.0 -26.55 162.6 ;
        RECT  -32.7 153.9 -32.1 154.5 ;
        RECT  -34.5 156.6 -33.9 157.2 ;
        RECT  -47.55 162.0 -46.95 162.6 ;
        RECT  -42.0 159.3 -41.4 159.9 ;
        RECT  -40.2 156.6 -39.6 157.2 ;
        RECT  -15.9 121.2 -15.3 121.8 ;
        RECT  -5.7 121.2 -5.1 121.8 ;
        RECT  -5.55 151.05 -4.95 151.65 ;
        RECT  -30.6 214.5 -30.0 215.1 ;
        RECT  -44.1 211.8 -43.5 212.4 ;
        RECT  -14.7 217.2 -14.1 217.8 ;
        RECT  -3.9 214.35 -3.3 214.95 ;
        RECT  -22.65 219.9 -22.05 220.5 ;
        RECT  -52.05 219.9 -51.45 220.5 ;
        RECT  -7.95 148.5 -7.35 149.1 ;
        RECT  -14.55 126.6 -13.95 127.2 ;
        RECT  -27.6 126.6 -27.0 127.2 ;
        RECT  -27.3 85.8 -26.7 86.4 ;
        RECT  -13.8 88.8 -13.2 89.4 ;
        RECT  -14.7 175.8 -14.1 176.4 ;
        RECT  -14.7 180.3 -14.1 180.9 ;
        RECT  0.3 219.9 0.9 220.5 ;
        RECT  1.5 219.9 2.1 220.5 ;
        Layer  metal2 ; 
        RECT  -7.5 219.6 0.0 220.5 ;
        RECT  95.1 0.0 104.1 459.3 ;
        RECT  119.4 0.0 120.3 459.3 ;
        RECT  116.7 0.0 117.6 459.3 ;
        RECT  114.0 0.0 114.9 459.3 ;
        RECT  111.3 0.0 112.2 459.3 ;
        RECT  108.6 0.0 109.5 459.3 ;
        RECT  105.9 0.0 106.8 459.3 ;
        RECT  90.6 39.0 91.5 196.5 ;
        RECT  87.9 39.0 88.8 196.5 ;
        RECT  85.2 39.0 86.1 196.5 ;
        RECT  82.5 39.0 83.4 196.5 ;
        RECT  127.05 435.3 127.95 439.8 ;
        RECT  130.05 435.3 130.95 439.8 ;
        RECT  137.25 435.3 138.15 439.8 ;
        RECT  140.25 435.3 141.15 439.8 ;
        RECT  147.45 435.3 148.35 439.8 ;
        RECT  150.45 435.3 151.35 439.8 ;
        RECT  114.0 200.1 114.9 448.2 ;
        RECT  133.65 435.3 134.55 438.0 ;
        RECT  143.85 435.3 144.75 438.0 ;
        RECT  154.05 435.3 154.95 438.0 ;
        RECT  123.0 200.1 123.9 438.0 ;
        RECT  88.5 229.05 95.1 229.95 ;
        RECT  88.5 258.45 95.1 259.35 ;
        RECT  88.5 287.85 95.1 288.75 ;
        RECT  88.5 317.25 95.1 318.15 ;
        RECT  88.5 346.65 95.1 347.55 ;
        RECT  88.5 376.05 95.1 376.95 ;
        RECT  88.5 405.45 95.1 406.35 ;
        RECT  88.5 434.85 95.1 435.75 ;
        RECT  123.3 204.3 125.7 214.8 ;
        RECT  126.9 201.3 128.1 214.8 ;
        RECT  129.9 201.3 131.1 214.8 ;
        RECT  125.4 200.1 128.1 201.3 ;
        RECT  129.6 200.1 131.1 201.3 ;
        RECT  133.5 200.1 134.7 214.8 ;
        RECT  123.3 214.8 125.7 225.3 ;
        RECT  126.9 214.8 128.1 228.3 ;
        RECT  129.9 214.8 131.1 228.3 ;
        RECT  125.4 228.3 128.1 229.5 ;
        RECT  129.6 228.3 131.1 229.5 ;
        RECT  133.5 214.8 134.7 229.5 ;
        RECT  123.3 233.7 125.7 244.2 ;
        RECT  126.9 230.7 128.1 244.2 ;
        RECT  129.9 230.7 131.1 244.2 ;
        RECT  125.4 229.5 128.1 230.7 ;
        RECT  129.6 229.5 131.1 230.7 ;
        RECT  133.5 229.5 134.7 244.2 ;
        RECT  123.3 244.2 125.7 254.7 ;
        RECT  126.9 244.2 128.1 257.7 ;
        RECT  129.9 244.2 131.1 257.7 ;
        RECT  125.4 257.7 128.1 258.9 ;
        RECT  129.6 257.7 131.1 258.9 ;
        RECT  133.5 244.2 134.7 258.9 ;
        RECT  123.3 263.1 125.7 273.6 ;
        RECT  126.9 260.1 128.1 273.6 ;
        RECT  129.9 260.1 131.1 273.6 ;
        RECT  125.4 258.9 128.1 260.1 ;
        RECT  129.6 258.9 131.1 260.1 ;
        RECT  133.5 258.9 134.7 273.6 ;
        RECT  123.3 273.6 125.7 284.1 ;
        RECT  126.9 273.6 128.1 287.1 ;
        RECT  129.9 273.6 131.1 287.1 ;
        RECT  125.4 287.1 128.1 288.3 ;
        RECT  129.6 287.1 131.1 288.3 ;
        RECT  133.5 273.6 134.7 288.3 ;
        RECT  123.3 292.5 125.7 303.0 ;
        RECT  126.9 289.5 128.1 303.0 ;
        RECT  129.9 289.5 131.1 303.0 ;
        RECT  125.4 288.3 128.1 289.5 ;
        RECT  129.6 288.3 131.1 289.5 ;
        RECT  133.5 288.3 134.7 303.0 ;
        RECT  123.3 303.0 125.7 313.5 ;
        RECT  126.9 303.0 128.1 316.5 ;
        RECT  129.9 303.0 131.1 316.5 ;
        RECT  125.4 316.5 128.1 317.7 ;
        RECT  129.6 316.5 131.1 317.7 ;
        RECT  133.5 303.0 134.7 317.7 ;
        RECT  123.3 321.9 125.7 332.4 ;
        RECT  126.9 318.9 128.1 332.4 ;
        RECT  129.9 318.9 131.1 332.4 ;
        RECT  125.4 317.7 128.1 318.9 ;
        RECT  129.6 317.7 131.1 318.9 ;
        RECT  133.5 317.7 134.7 332.4 ;
        RECT  123.3 332.4 125.7 342.9 ;
        RECT  126.9 332.4 128.1 345.9 ;
        RECT  129.9 332.4 131.1 345.9 ;
        RECT  125.4 345.9 128.1 347.1 ;
        RECT  129.6 345.9 131.1 347.1 ;
        RECT  133.5 332.4 134.7 347.1 ;
        RECT  123.3 351.3 125.7 361.8 ;
        RECT  126.9 348.3 128.1 361.8 ;
        RECT  129.9 348.3 131.1 361.8 ;
        RECT  125.4 347.1 128.1 348.3 ;
        RECT  129.6 347.1 131.1 348.3 ;
        RECT  133.5 347.1 134.7 361.8 ;
        RECT  123.3 361.8 125.7 372.3 ;
        RECT  126.9 361.8 128.1 375.3 ;
        RECT  129.9 361.8 131.1 375.3 ;
        RECT  125.4 375.3 128.1 376.5 ;
        RECT  129.6 375.3 131.1 376.5 ;
        RECT  133.5 361.8 134.7 376.5 ;
        RECT  123.3 380.7 125.7 391.2 ;
        RECT  126.9 377.7 128.1 391.2 ;
        RECT  129.9 377.7 131.1 391.2 ;
        RECT  125.4 376.5 128.1 377.7 ;
        RECT  129.6 376.5 131.1 377.7 ;
        RECT  133.5 376.5 134.7 391.2 ;
        RECT  123.3 391.2 125.7 401.7 ;
        RECT  126.9 391.2 128.1 404.7 ;
        RECT  129.9 391.2 131.1 404.7 ;
        RECT  125.4 404.7 128.1 405.9 ;
        RECT  129.6 404.7 131.1 405.9 ;
        RECT  133.5 391.2 134.7 405.9 ;
        RECT  123.3 410.1 125.7 420.6 ;
        RECT  126.9 407.1 128.1 420.6 ;
        RECT  129.9 407.1 131.1 420.6 ;
        RECT  125.4 405.9 128.1 407.1 ;
        RECT  129.6 405.9 131.1 407.1 ;
        RECT  133.5 405.9 134.7 420.6 ;
        RECT  123.3 420.6 125.7 431.1 ;
        RECT  126.9 420.6 128.1 434.1 ;
        RECT  129.9 420.6 131.1 434.1 ;
        RECT  125.4 434.1 128.1 435.3 ;
        RECT  129.6 434.1 131.1 435.3 ;
        RECT  133.5 420.6 134.7 435.3 ;
        RECT  133.5 204.3 135.9 214.8 ;
        RECT  137.1 201.3 138.3 214.8 ;
        RECT  140.1 201.3 141.3 214.8 ;
        RECT  135.6 200.1 138.3 201.3 ;
        RECT  139.8 200.1 141.3 201.3 ;
        RECT  143.7 200.1 144.9 214.8 ;
        RECT  133.5 214.8 135.9 225.3 ;
        RECT  137.1 214.8 138.3 228.3 ;
        RECT  140.1 214.8 141.3 228.3 ;
        RECT  135.6 228.3 138.3 229.5 ;
        RECT  139.8 228.3 141.3 229.5 ;
        RECT  143.7 214.8 144.9 229.5 ;
        RECT  133.5 233.7 135.9 244.2 ;
        RECT  137.1 230.7 138.3 244.2 ;
        RECT  140.1 230.7 141.3 244.2 ;
        RECT  135.6 229.5 138.3 230.7 ;
        RECT  139.8 229.5 141.3 230.7 ;
        RECT  143.7 229.5 144.9 244.2 ;
        RECT  133.5 244.2 135.9 254.7 ;
        RECT  137.1 244.2 138.3 257.7 ;
        RECT  140.1 244.2 141.3 257.7 ;
        RECT  135.6 257.7 138.3 258.9 ;
        RECT  139.8 257.7 141.3 258.9 ;
        RECT  143.7 244.2 144.9 258.9 ;
        RECT  133.5 263.1 135.9 273.6 ;
        RECT  137.1 260.1 138.3 273.6 ;
        RECT  140.1 260.1 141.3 273.6 ;
        RECT  135.6 258.9 138.3 260.1 ;
        RECT  139.8 258.9 141.3 260.1 ;
        RECT  143.7 258.9 144.9 273.6 ;
        RECT  133.5 273.6 135.9 284.1 ;
        RECT  137.1 273.6 138.3 287.1 ;
        RECT  140.1 273.6 141.3 287.1 ;
        RECT  135.6 287.1 138.3 288.3 ;
        RECT  139.8 287.1 141.3 288.3 ;
        RECT  143.7 273.6 144.9 288.3 ;
        RECT  133.5 292.5 135.9 303.0 ;
        RECT  137.1 289.5 138.3 303.0 ;
        RECT  140.1 289.5 141.3 303.0 ;
        RECT  135.6 288.3 138.3 289.5 ;
        RECT  139.8 288.3 141.3 289.5 ;
        RECT  143.7 288.3 144.9 303.0 ;
        RECT  133.5 303.0 135.9 313.5 ;
        RECT  137.1 303.0 138.3 316.5 ;
        RECT  140.1 303.0 141.3 316.5 ;
        RECT  135.6 316.5 138.3 317.7 ;
        RECT  139.8 316.5 141.3 317.7 ;
        RECT  143.7 303.0 144.9 317.7 ;
        RECT  133.5 321.9 135.9 332.4 ;
        RECT  137.1 318.9 138.3 332.4 ;
        RECT  140.1 318.9 141.3 332.4 ;
        RECT  135.6 317.7 138.3 318.9 ;
        RECT  139.8 317.7 141.3 318.9 ;
        RECT  143.7 317.7 144.9 332.4 ;
        RECT  133.5 332.4 135.9 342.9 ;
        RECT  137.1 332.4 138.3 345.9 ;
        RECT  140.1 332.4 141.3 345.9 ;
        RECT  135.6 345.9 138.3 347.1 ;
        RECT  139.8 345.9 141.3 347.1 ;
        RECT  143.7 332.4 144.9 347.1 ;
        RECT  133.5 351.3 135.9 361.8 ;
        RECT  137.1 348.3 138.3 361.8 ;
        RECT  140.1 348.3 141.3 361.8 ;
        RECT  135.6 347.1 138.3 348.3 ;
        RECT  139.8 347.1 141.3 348.3 ;
        RECT  143.7 347.1 144.9 361.8 ;
        RECT  133.5 361.8 135.9 372.3 ;
        RECT  137.1 361.8 138.3 375.3 ;
        RECT  140.1 361.8 141.3 375.3 ;
        RECT  135.6 375.3 138.3 376.5 ;
        RECT  139.8 375.3 141.3 376.5 ;
        RECT  143.7 361.8 144.9 376.5 ;
        RECT  133.5 380.7 135.9 391.2 ;
        RECT  137.1 377.7 138.3 391.2 ;
        RECT  140.1 377.7 141.3 391.2 ;
        RECT  135.6 376.5 138.3 377.7 ;
        RECT  139.8 376.5 141.3 377.7 ;
        RECT  143.7 376.5 144.9 391.2 ;
        RECT  133.5 391.2 135.9 401.7 ;
        RECT  137.1 391.2 138.3 404.7 ;
        RECT  140.1 391.2 141.3 404.7 ;
        RECT  135.6 404.7 138.3 405.9 ;
        RECT  139.8 404.7 141.3 405.9 ;
        RECT  143.7 391.2 144.9 405.9 ;
        RECT  133.5 410.1 135.9 420.6 ;
        RECT  137.1 407.1 138.3 420.6 ;
        RECT  140.1 407.1 141.3 420.6 ;
        RECT  135.6 405.9 138.3 407.1 ;
        RECT  139.8 405.9 141.3 407.1 ;
        RECT  143.7 405.9 144.9 420.6 ;
        RECT  133.5 420.6 135.9 431.1 ;
        RECT  137.1 420.6 138.3 434.1 ;
        RECT  140.1 420.6 141.3 434.1 ;
        RECT  135.6 434.1 138.3 435.3 ;
        RECT  139.8 434.1 141.3 435.3 ;
        RECT  143.7 420.6 144.9 435.3 ;
        RECT  143.7 204.3 146.1 214.8 ;
        RECT  147.3 201.3 148.5 214.8 ;
        RECT  150.3 201.3 151.5 214.8 ;
        RECT  145.8 200.1 148.5 201.3 ;
        RECT  150.0 200.1 151.5 201.3 ;
        RECT  153.9 200.1 155.1 214.8 ;
        RECT  143.7 214.8 146.1 225.3 ;
        RECT  147.3 214.8 148.5 228.3 ;
        RECT  150.3 214.8 151.5 228.3 ;
        RECT  145.8 228.3 148.5 229.5 ;
        RECT  150.0 228.3 151.5 229.5 ;
        RECT  153.9 214.8 155.1 229.5 ;
        RECT  143.7 233.7 146.1 244.2 ;
        RECT  147.3 230.7 148.5 244.2 ;
        RECT  150.3 230.7 151.5 244.2 ;
        RECT  145.8 229.5 148.5 230.7 ;
        RECT  150.0 229.5 151.5 230.7 ;
        RECT  153.9 229.5 155.1 244.2 ;
        RECT  143.7 244.2 146.1 254.7 ;
        RECT  147.3 244.2 148.5 257.7 ;
        RECT  150.3 244.2 151.5 257.7 ;
        RECT  145.8 257.7 148.5 258.9 ;
        RECT  150.0 257.7 151.5 258.9 ;
        RECT  153.9 244.2 155.1 258.9 ;
        RECT  143.7 263.1 146.1 273.6 ;
        RECT  147.3 260.1 148.5 273.6 ;
        RECT  150.3 260.1 151.5 273.6 ;
        RECT  145.8 258.9 148.5 260.1 ;
        RECT  150.0 258.9 151.5 260.1 ;
        RECT  153.9 258.9 155.1 273.6 ;
        RECT  143.7 273.6 146.1 284.1 ;
        RECT  147.3 273.6 148.5 287.1 ;
        RECT  150.3 273.6 151.5 287.1 ;
        RECT  145.8 287.1 148.5 288.3 ;
        RECT  150.0 287.1 151.5 288.3 ;
        RECT  153.9 273.6 155.1 288.3 ;
        RECT  143.7 292.5 146.1 303.0 ;
        RECT  147.3 289.5 148.5 303.0 ;
        RECT  150.3 289.5 151.5 303.0 ;
        RECT  145.8 288.3 148.5 289.5 ;
        RECT  150.0 288.3 151.5 289.5 ;
        RECT  153.9 288.3 155.1 303.0 ;
        RECT  143.7 303.0 146.1 313.5 ;
        RECT  147.3 303.0 148.5 316.5 ;
        RECT  150.3 303.0 151.5 316.5 ;
        RECT  145.8 316.5 148.5 317.7 ;
        RECT  150.0 316.5 151.5 317.7 ;
        RECT  153.9 303.0 155.1 317.7 ;
        RECT  143.7 321.9 146.1 332.4 ;
        RECT  147.3 318.9 148.5 332.4 ;
        RECT  150.3 318.9 151.5 332.4 ;
        RECT  145.8 317.7 148.5 318.9 ;
        RECT  150.0 317.7 151.5 318.9 ;
        RECT  153.9 317.7 155.1 332.4 ;
        RECT  143.7 332.4 146.1 342.9 ;
        RECT  147.3 332.4 148.5 345.9 ;
        RECT  150.3 332.4 151.5 345.9 ;
        RECT  145.8 345.9 148.5 347.1 ;
        RECT  150.0 345.9 151.5 347.1 ;
        RECT  153.9 332.4 155.1 347.1 ;
        RECT  143.7 351.3 146.1 361.8 ;
        RECT  147.3 348.3 148.5 361.8 ;
        RECT  150.3 348.3 151.5 361.8 ;
        RECT  145.8 347.1 148.5 348.3 ;
        RECT  150.0 347.1 151.5 348.3 ;
        RECT  153.9 347.1 155.1 361.8 ;
        RECT  143.7 361.8 146.1 372.3 ;
        RECT  147.3 361.8 148.5 375.3 ;
        RECT  150.3 361.8 151.5 375.3 ;
        RECT  145.8 375.3 148.5 376.5 ;
        RECT  150.0 375.3 151.5 376.5 ;
        RECT  153.9 361.8 155.1 376.5 ;
        RECT  143.7 380.7 146.1 391.2 ;
        RECT  147.3 377.7 148.5 391.2 ;
        RECT  150.3 377.7 151.5 391.2 ;
        RECT  145.8 376.5 148.5 377.7 ;
        RECT  150.0 376.5 151.5 377.7 ;
        RECT  153.9 376.5 155.1 391.2 ;
        RECT  143.7 391.2 146.1 401.7 ;
        RECT  147.3 391.2 148.5 404.7 ;
        RECT  150.3 391.2 151.5 404.7 ;
        RECT  145.8 404.7 148.5 405.9 ;
        RECT  150.0 404.7 151.5 405.9 ;
        RECT  153.9 391.2 155.1 405.9 ;
        RECT  143.7 410.1 146.1 420.6 ;
        RECT  147.3 407.1 148.5 420.6 ;
        RECT  150.3 407.1 151.5 420.6 ;
        RECT  145.8 405.9 148.5 407.1 ;
        RECT  150.0 405.9 151.5 407.1 ;
        RECT  153.9 405.9 155.1 420.6 ;
        RECT  143.7 420.6 146.1 431.1 ;
        RECT  147.3 420.6 148.5 434.1 ;
        RECT  150.3 420.6 151.5 434.1 ;
        RECT  145.8 434.1 148.5 435.3 ;
        RECT  150.0 434.1 151.5 435.3 ;
        RECT  153.9 420.6 155.1 435.3 ;
        RECT  127.05 439.8 127.95 459.3 ;
        RECT  130.05 439.8 130.95 459.3 ;
        RECT  127.35 450.9 127.5 452.1 ;
        RECT  130.05 450.9 131.7 452.1 ;
        RECT  127.35 442.5 127.5 443.7 ;
        RECT  129.3 442.5 130.05 443.7 ;
        RECT  126.9 450.9 128.1 452.1 ;
        RECT  131.7 450.9 132.9 452.1 ;
        RECT  126.9 442.5 128.1 443.7 ;
        RECT  129.3 442.5 130.5 443.7 ;
        RECT  137.25 439.8 138.15 459.3 ;
        RECT  140.25 439.8 141.15 459.3 ;
        RECT  137.55 450.9 137.7 452.1 ;
        RECT  140.25 450.9 141.9 452.1 ;
        RECT  137.55 442.5 137.7 443.7 ;
        RECT  139.5 442.5 140.25 443.7 ;
        RECT  137.1 450.9 138.3 452.1 ;
        RECT  141.9 450.9 143.1 452.1 ;
        RECT  137.1 442.5 138.3 443.7 ;
        RECT  139.5 442.5 140.7 443.7 ;
        RECT  147.45 439.8 148.35 459.3 ;
        RECT  150.45 439.8 151.35 459.3 ;
        RECT  147.75 450.9 147.9 452.1 ;
        RECT  150.45 450.9 152.1 452.1 ;
        RECT  147.75 442.5 147.9 443.7 ;
        RECT  149.7 442.5 150.45 443.7 ;
        RECT  147.3 450.9 148.5 452.1 ;
        RECT  152.1 450.9 153.3 452.1 ;
        RECT  147.3 442.5 148.5 443.7 ;
        RECT  149.7 442.5 150.9 443.7 ;
        RECT  126.9 165.6 128.1 200.1 ;
        RECT  129.9 165.6 131.1 200.1 ;
        RECT  133.5 192.6 134.7 200.1 ;
        RECT  126.9 164.4 129.0 165.6 ;
        RECT  129.9 164.4 131.7 165.6 ;
        RECT  124.8 151.2 126.0 155.7 ;
        RECT  126.9 151.2 128.1 164.4 ;
        RECT  129.9 151.2 131.1 164.4 ;
        RECT  137.1 165.6 138.3 200.1 ;
        RECT  140.1 165.6 141.3 200.1 ;
        RECT  143.7 192.6 144.9 200.1 ;
        RECT  137.1 164.4 139.2 165.6 ;
        RECT  140.1 164.4 141.9 165.6 ;
        RECT  135.0 151.2 136.2 155.7 ;
        RECT  137.1 151.2 138.3 164.4 ;
        RECT  140.1 151.2 141.3 164.4 ;
        RECT  147.3 165.6 148.5 200.1 ;
        RECT  150.3 165.6 151.5 200.1 ;
        RECT  153.9 192.6 155.1 200.1 ;
        RECT  147.3 164.4 149.4 165.6 ;
        RECT  150.3 164.4 152.1 165.6 ;
        RECT  145.2 151.2 146.4 155.7 ;
        RECT  147.3 151.2 148.5 164.4 ;
        RECT  150.3 151.2 151.5 164.4 ;
        RECT  126.9 149.1 128.1 151.2 ;
        RECT  125.4 147.9 128.1 149.1 ;
        RECT  129.9 143.7 131.1 151.2 ;
        RECT  133.5 138.9 134.7 149.4 ;
        RECT  127.2 137.7 134.7 138.9 ;
        RECT  126.3 99.9 127.5 127.2 ;
        RECT  133.5 116.4 134.7 137.7 ;
        RECT  132.9 115.2 134.7 116.4 ;
        RECT  133.5 112.2 134.7 115.2 ;
        RECT  129.6 111.0 134.7 112.2 ;
        RECT  129.6 109.8 130.8 111.0 ;
        RECT  127.5 93.6 129.9 94.8 ;
        RECT  128.4 90.9 129.6 93.6 ;
        RECT  133.5 90.9 134.7 111.0 ;
        RECT  137.1 149.1 138.3 151.2 ;
        RECT  135.6 147.9 138.3 149.1 ;
        RECT  140.1 143.7 141.3 151.2 ;
        RECT  143.7 138.9 144.9 149.4 ;
        RECT  137.4 137.7 144.9 138.9 ;
        RECT  136.5 99.9 137.7 127.2 ;
        RECT  143.7 116.4 144.9 137.7 ;
        RECT  143.1 115.2 144.9 116.4 ;
        RECT  143.7 112.2 144.9 115.2 ;
        RECT  139.8 111.0 144.9 112.2 ;
        RECT  139.8 109.8 141.0 111.0 ;
        RECT  137.7 93.6 140.1 94.8 ;
        RECT  138.6 90.9 139.8 93.6 ;
        RECT  143.7 90.9 144.9 111.0 ;
        RECT  147.3 149.1 148.5 151.2 ;
        RECT  145.8 147.9 148.5 149.1 ;
        RECT  150.3 143.7 151.5 151.2 ;
        RECT  153.9 138.9 155.1 149.4 ;
        RECT  147.6 137.7 155.1 138.9 ;
        RECT  146.7 99.9 147.9 127.2 ;
        RECT  153.9 116.4 155.1 137.7 ;
        RECT  153.3 115.2 155.1 116.4 ;
        RECT  153.9 112.2 155.1 115.2 ;
        RECT  150.0 111.0 155.1 112.2 ;
        RECT  150.0 109.8 151.2 111.0 ;
        RECT  147.9 93.6 150.3 94.8 ;
        RECT  148.8 90.9 150.0 93.6 ;
        RECT  153.9 90.9 155.1 111.0 ;
        RECT  125.7 86.4 126.9 90.9 ;
        RECT  128.4 89.7 129.6 90.9 ;
        RECT  128.4 88.5 131.1 89.7 ;
        RECT  125.7 85.2 128.7 86.4 ;
        RECT  125.7 75.6 126.6 85.2 ;
        RECT  129.9 80.7 131.1 88.5 ;
        RECT  129.0 77.4 132.0 78.6 ;
        RECT  125.7 74.4 126.9 75.6 ;
        RECT  129.0 75.3 130.2 76.5 ;
        RECT  129.3 73.8 130.2 75.3 ;
        RECT  127.8 72.9 130.2 73.8 ;
        RECT  127.8 66.6 128.7 72.9 ;
        RECT  131.1 72.0 132.0 77.4 ;
        RECT  129.9 70.8 132.0 72.0 ;
        RECT  129.9 68.4 132.0 69.6 ;
        RECT  127.5 65.4 128.7 66.6 ;
        RECT  125.4 60.9 126.9 62.1 ;
        RECT  125.4 49.2 126.3 60.9 ;
        RECT  128.4 58.8 129.6 63.3 ;
        RECT  127.2 57.9 129.6 58.8 ;
        RECT  127.2 51.0 128.1 57.9 ;
        RECT  131.1 56.4 132.0 68.4 ;
        RECT  129.9 55.2 132.0 56.4 ;
        RECT  129.0 51.9 132.0 53.1 ;
        RECT  127.2 50.1 128.7 51.0 ;
        RECT  125.4 48.0 126.9 49.2 ;
        RECT  127.8 48.9 130.2 50.1 ;
        RECT  127.8 40.2 128.7 48.9 ;
        RECT  131.1 45.6 132.0 51.9 ;
        RECT  129.9 44.4 132.0 45.6 ;
        RECT  129.9 42.0 132.0 43.2 ;
        RECT  127.5 39.0 128.7 40.2 ;
        RECT  131.1 33.3 132.0 42.0 ;
        RECT  128.4 32.1 132.0 33.3 ;
        RECT  128.4 30.9 129.6 32.1 ;
        RECT  133.5 30.9 134.7 90.9 ;
        RECT  141.3 86.4 142.5 90.9 ;
        RECT  138.6 89.7 139.8 90.9 ;
        RECT  137.1 88.5 139.8 89.7 ;
        RECT  139.5 85.2 142.5 86.4 ;
        RECT  141.6 75.6 142.5 85.2 ;
        RECT  137.1 80.7 138.3 88.5 ;
        RECT  136.2 77.4 139.2 78.6 ;
        RECT  141.3 74.4 142.5 75.6 ;
        RECT  138.0 75.3 139.2 76.5 ;
        RECT  138.0 73.8 138.9 75.3 ;
        RECT  138.0 72.9 140.4 73.8 ;
        RECT  139.5 66.6 140.4 72.9 ;
        RECT  136.2 72.0 137.1 77.4 ;
        RECT  136.2 70.8 138.3 72.0 ;
        RECT  136.2 68.4 138.3 69.6 ;
        RECT  139.5 65.4 140.7 66.6 ;
        RECT  141.3 60.9 142.8 62.1 ;
        RECT  141.9 49.2 142.8 60.9 ;
        RECT  138.6 58.8 139.8 63.3 ;
        RECT  138.6 57.9 141.0 58.8 ;
        RECT  140.1 51.0 141.0 57.9 ;
        RECT  136.2 56.4 137.1 68.4 ;
        RECT  136.2 55.2 138.3 56.4 ;
        RECT  136.2 51.9 139.2 53.1 ;
        RECT  139.5 50.1 141.0 51.0 ;
        RECT  141.3 48.0 142.8 49.2 ;
        RECT  138.0 48.9 140.4 50.1 ;
        RECT  139.5 40.2 140.4 48.9 ;
        RECT  136.2 45.6 137.1 51.9 ;
        RECT  136.2 44.4 138.3 45.6 ;
        RECT  136.2 42.0 138.3 43.2 ;
        RECT  139.5 39.0 140.7 40.2 ;
        RECT  136.2 33.3 137.1 42.0 ;
        RECT  136.2 32.1 139.8 33.3 ;
        RECT  138.6 30.9 139.8 32.1 ;
        RECT  133.5 30.9 134.7 90.9 ;
        RECT  146.1 86.4 147.3 90.9 ;
        RECT  148.8 89.7 150.0 90.9 ;
        RECT  148.8 88.5 151.5 89.7 ;
        RECT  146.1 85.2 149.1 86.4 ;
        RECT  146.1 75.6 147.0 85.2 ;
        RECT  150.3 80.7 151.5 88.5 ;
        RECT  149.4 77.4 152.4 78.6 ;
        RECT  146.1 74.4 147.3 75.6 ;
        RECT  149.4 75.3 150.6 76.5 ;
        RECT  149.7 73.8 150.6 75.3 ;
        RECT  148.2 72.9 150.6 73.8 ;
        RECT  148.2 66.6 149.1 72.9 ;
        RECT  151.5 72.0 152.4 77.4 ;
        RECT  150.3 70.8 152.4 72.0 ;
        RECT  150.3 68.4 152.4 69.6 ;
        RECT  147.9 65.4 149.1 66.6 ;
        RECT  145.8 60.9 147.3 62.1 ;
        RECT  145.8 49.2 146.7 60.9 ;
        RECT  148.8 58.8 150.0 63.3 ;
        RECT  147.6 57.9 150.0 58.8 ;
        RECT  147.6 51.0 148.5 57.9 ;
        RECT  151.5 56.4 152.4 68.4 ;
        RECT  150.3 55.2 152.4 56.4 ;
        RECT  149.4 51.9 152.4 53.1 ;
        RECT  147.6 50.1 149.1 51.0 ;
        RECT  145.8 48.0 147.3 49.2 ;
        RECT  148.2 48.9 150.6 50.1 ;
        RECT  148.2 40.2 149.1 48.9 ;
        RECT  151.5 45.6 152.4 51.9 ;
        RECT  150.3 44.4 152.4 45.6 ;
        RECT  150.3 42.0 152.4 43.2 ;
        RECT  147.9 39.0 149.1 40.2 ;
        RECT  151.5 33.3 152.4 42.0 ;
        RECT  148.8 32.1 152.4 33.3 ;
        RECT  148.8 30.9 150.0 32.1 ;
        RECT  153.9 30.9 155.1 90.9 ;
        RECT  128.4 45.9 129.6 52.8 ;
        RECT  126.6 44.7 129.6 45.9 ;
        RECT  128.4 41.1 132.6 42.3 ;
        RECT  128.4 33.6 129.6 41.1 ;
        RECT  128.4 32.4 129.9 33.6 ;
        RECT  128.4 30.9 129.6 32.4 ;
        RECT  133.5 30.9 134.7 52.8 ;
        RECT  138.6 45.9 139.8 52.8 ;
        RECT  138.6 44.7 141.6 45.9 ;
        RECT  135.6 41.1 139.8 42.3 ;
        RECT  138.6 33.6 139.8 41.1 ;
        RECT  138.3 32.4 139.8 33.6 ;
        RECT  138.6 30.9 139.8 32.4 ;
        RECT  133.5 30.9 134.7 52.8 ;
        RECT  148.8 45.9 150.0 52.8 ;
        RECT  147.0 44.7 150.0 45.9 ;
        RECT  148.8 41.1 153.0 42.3 ;
        RECT  148.8 33.6 150.0 41.1 ;
        RECT  148.8 32.4 150.3 33.6 ;
        RECT  148.8 30.9 150.0 32.4 ;
        RECT  153.9 30.9 155.1 52.8 ;
        RECT  27.3 82.5 28.2 435.3 ;
        RECT  25.2 82.5 26.1 435.3 ;
        RECT  23.1 82.5 24.0 435.3 ;
        RECT  21.0 82.5 21.9 435.3 ;
        RECT  18.9 82.5 19.8 435.3 ;
        RECT  16.8 82.5 17.7 435.3 ;
        RECT  14.7 82.5 15.6 435.3 ;
        RECT  12.6 82.5 13.5 435.3 ;
        RECT  77.7 82.5 78.6 138.6 ;
        RECT  75.6 82.5 76.5 138.6 ;
        RECT  62.7 82.5 63.6 138.6 ;
        RECT  60.6 82.5 61.5 138.6 ;
        RECT  58.5 82.5 59.4 138.6 ;
        RECT  56.4 82.5 57.3 138.6 ;
        RECT  54.3 82.5 55.2 138.6 ;
        RECT  52.2 82.5 53.1 138.6 ;
        RECT  58.2 92.85 59.4 94.05 ;
        RECT  77.4 87.6 78.6 88.8 ;
        RECT  56.1 98.25 57.3 99.45 ;
        RECT  75.3 103.5 76.5 104.7 ;
        RECT  58.2 90.0 59.4 91.2 ;
        RECT  56.1 86.7 57.3 87.9 ;
        RECT  54.0 101.1 55.2 102.3 ;
        RECT  56.1 104.4 57.3 105.6 ;
        RECT  58.2 119.4 59.4 120.6 ;
        RECT  51.9 116.1 53.1 117.3 ;
        RECT  54.0 130.5 55.2 131.7 ;
        RECT  77.4 130.5 78.6 131.7 ;
        RECT  51.9 133.8 53.1 135.0 ;
        RECT  75.3 133.8 76.5 135.0 ;
        RECT  60.3 80.85 61.5 82.05 ;
        RECT  62.4 95.55 63.6 96.75 ;
        RECT  60.3 110.25 61.5 111.45 ;
        RECT  62.4 124.95 63.6 126.15 ;
        RECT  60.3 137.4 61.5 138.6 ;
        RECT  77.7 141.3 78.6 197.4 ;
        RECT  75.6 141.3 76.5 197.4 ;
        RECT  62.7 141.3 63.6 197.4 ;
        RECT  60.6 141.3 61.5 197.4 ;
        RECT  58.5 141.3 59.4 197.4 ;
        RECT  56.4 141.3 57.3 197.4 ;
        RECT  54.3 141.3 55.2 197.4 ;
        RECT  52.2 141.3 53.1 197.4 ;
        RECT  58.2 151.65 59.4 152.85 ;
        RECT  77.4 146.4 78.6 147.6 ;
        RECT  56.1 157.05 57.3 158.25 ;
        RECT  75.3 162.3 76.5 163.5 ;
        RECT  58.2 148.8 59.4 150.0 ;
        RECT  56.1 145.5 57.3 146.7 ;
        RECT  54.0 159.9 55.2 161.1 ;
        RECT  56.1 163.2 57.3 164.4 ;
        RECT  58.2 178.2 59.4 179.4 ;
        RECT  51.9 174.9 53.1 176.1 ;
        RECT  54.0 189.3 55.2 190.5 ;
        RECT  77.4 189.3 78.6 190.5 ;
        RECT  51.9 192.6 53.1 193.8 ;
        RECT  75.3 192.6 76.5 193.8 ;
        RECT  60.3 139.65 61.5 140.85 ;
        RECT  62.4 154.35 63.6 155.55 ;
        RECT  60.3 169.05 61.5 170.25 ;
        RECT  62.4 183.75 63.6 184.95 ;
        RECT  60.3 196.2 61.5 197.4 ;
        RECT  12.6 88.8 13.8 90.0 ;
        RECT  14.7 104.7 15.9 105.9 ;
        RECT  16.8 118.2 18.0 119.4 ;
        RECT  18.9 134.1 20.1 135.3 ;
        RECT  21.0 147.6 22.2 148.8 ;
        RECT  23.1 163.5 24.3 164.7 ;
        RECT  25.2 177.0 26.4 178.2 ;
        RECT  27.3 192.9 28.5 194.1 ;
        RECT  12.6 208.8 13.8 210.0 ;
        RECT  21.0 205.5 22.2 206.7 ;
        RECT  12.6 219.9 13.8 221.1 ;
        RECT  23.1 223.2 24.3 224.4 ;
        RECT  12.6 238.2 13.8 239.4 ;
        RECT  25.2 234.9 26.4 236.1 ;
        RECT  12.6 249.3 13.8 250.5 ;
        RECT  27.3 252.6 28.5 253.8 ;
        RECT  14.7 267.6 15.9 268.8 ;
        RECT  21.0 264.3 22.2 265.5 ;
        RECT  14.7 278.7 15.9 279.9 ;
        RECT  23.1 282.0 24.3 283.2 ;
        RECT  14.7 297.0 15.9 298.2 ;
        RECT  25.2 293.7 26.4 294.9 ;
        RECT  14.7 308.1 15.9 309.3 ;
        RECT  27.3 311.4 28.5 312.6 ;
        RECT  16.8 326.4 18.0 327.6 ;
        RECT  21.0 323.1 22.2 324.3 ;
        RECT  16.8 337.5 18.0 338.7 ;
        RECT  23.1 340.8 24.3 342.0 ;
        RECT  16.8 355.8 18.0 357.0 ;
        RECT  25.2 352.5 26.4 353.7 ;
        RECT  16.8 366.9 18.0 368.1 ;
        RECT  27.3 370.2 28.5 371.4 ;
        RECT  18.9 385.2 20.1 386.4 ;
        RECT  21.0 381.9 22.2 383.1 ;
        RECT  18.9 396.3 20.1 397.5 ;
        RECT  23.1 399.6 24.3 400.8 ;
        RECT  18.9 414.6 20.1 415.8 ;
        RECT  25.2 411.3 26.4 412.5 ;
        RECT  18.9 425.7 20.1 426.9 ;
        RECT  27.3 429.0 28.5 430.2 ;
        RECT  51.0 214.35 57.3 215.25 ;
        RECT  51.0 208.8 66.9 209.7 ;
        RECT  51.0 229.05 57.3 229.95 ;
        RECT  51.0 219.9 66.9 220.8 ;
        RECT  51.0 243.75 57.3 244.65 ;
        RECT  51.0 238.2 66.9 239.1 ;
        RECT  51.0 258.45 57.3 259.35 ;
        RECT  51.0 249.3 66.9 250.2 ;
        RECT  51.0 273.15 57.3 274.05 ;
        RECT  51.0 267.6 66.9 268.5 ;
        RECT  51.0 287.85 57.3 288.75 ;
        RECT  51.0 278.7 66.9 279.6 ;
        RECT  51.0 302.55 57.3 303.45 ;
        RECT  51.0 297.0 66.9 297.9 ;
        RECT  51.0 317.25 57.3 318.15 ;
        RECT  51.0 308.1 66.9 309.0 ;
        RECT  51.0 331.95 57.3 332.85 ;
        RECT  51.0 326.4 66.9 327.3 ;
        RECT  51.0 346.65 57.3 347.55 ;
        RECT  51.0 337.5 66.9 338.4 ;
        RECT  51.0 361.35 57.3 362.25 ;
        RECT  51.0 355.8 66.9 356.7 ;
        RECT  51.0 376.05 57.3 376.95 ;
        RECT  51.0 366.9 66.9 367.8 ;
        RECT  51.0 390.75 57.3 391.65 ;
        RECT  51.0 385.2 66.9 386.1 ;
        RECT  51.0 405.45 57.3 406.35 ;
        RECT  51.0 396.3 66.9 397.2 ;
        RECT  51.0 420.15 57.3 421.05 ;
        RECT  51.0 414.6 66.9 415.5 ;
        RECT  51.0 434.85 57.3 435.75 ;
        RECT  51.0 425.7 66.9 426.6 ;
        RECT  50.7 214.35 51.9 215.55 ;
        RECT  57.0 214.35 58.2 215.55 ;
        RECT  66.9 208.8 68.1 210.0 ;
        RECT  51.0 208.8 52.2 210.0 ;
        RECT  50.7 229.05 51.9 230.25 ;
        RECT  57.0 229.05 58.2 230.25 ;
        RECT  66.9 219.6 68.1 220.8 ;
        RECT  51.0 219.6 52.2 220.8 ;
        RECT  50.7 243.75 51.9 244.95 ;
        RECT  57.0 243.75 58.2 244.95 ;
        RECT  66.9 238.2 68.1 239.4 ;
        RECT  51.0 238.2 52.2 239.4 ;
        RECT  50.7 258.45 51.9 259.65 ;
        RECT  57.0 258.45 58.2 259.65 ;
        RECT  66.9 249.0 68.1 250.2 ;
        RECT  51.0 249.0 52.2 250.2 ;
        RECT  50.7 273.15 51.9 274.35 ;
        RECT  57.0 273.15 58.2 274.35 ;
        RECT  66.9 267.6 68.1 268.8 ;
        RECT  51.0 267.6 52.2 268.8 ;
        RECT  50.7 287.85 51.9 289.05 ;
        RECT  57.0 287.85 58.2 289.05 ;
        RECT  66.9 278.4 68.1 279.6 ;
        RECT  51.0 278.4 52.2 279.6 ;
        RECT  50.7 302.55 51.9 303.75 ;
        RECT  57.0 302.55 58.2 303.75 ;
        RECT  66.9 297.0 68.1 298.2 ;
        RECT  51.0 297.0 52.2 298.2 ;
        RECT  50.7 317.25 51.9 318.45 ;
        RECT  57.0 317.25 58.2 318.45 ;
        RECT  66.9 307.8 68.1 309.0 ;
        RECT  51.0 307.8 52.2 309.0 ;
        RECT  50.7 331.95 51.9 333.15 ;
        RECT  57.0 331.95 58.2 333.15 ;
        RECT  66.9 326.4 68.1 327.6 ;
        RECT  51.0 326.4 52.2 327.6 ;
        RECT  50.7 346.65 51.9 347.85 ;
        RECT  57.0 346.65 58.2 347.85 ;
        RECT  66.9 337.2 68.1 338.4 ;
        RECT  51.0 337.2 52.2 338.4 ;
        RECT  50.7 361.35 51.9 362.55 ;
        RECT  57.0 361.35 58.2 362.55 ;
        RECT  66.9 355.8 68.1 357.0 ;
        RECT  51.0 355.8 52.2 357.0 ;
        RECT  50.7 376.05 51.9 377.25 ;
        RECT  57.0 376.05 58.2 377.25 ;
        RECT  66.9 366.6 68.1 367.8 ;
        RECT  51.0 366.6 52.2 367.8 ;
        RECT  50.7 390.75 51.9 391.95 ;
        RECT  57.0 390.75 58.2 391.95 ;
        RECT  66.9 385.2 68.1 386.4 ;
        RECT  51.0 385.2 52.2 386.4 ;
        RECT  50.7 405.45 51.9 406.65 ;
        RECT  57.0 405.45 58.2 406.65 ;
        RECT  66.9 396.0 68.1 397.2 ;
        RECT  51.0 396.0 52.2 397.2 ;
        RECT  50.7 420.15 51.9 421.35 ;
        RECT  57.0 420.15 58.2 421.35 ;
        RECT  66.9 414.6 68.1 415.8 ;
        RECT  51.0 414.6 52.2 415.8 ;
        RECT  50.7 434.85 51.9 436.05 ;
        RECT  57.0 434.85 58.2 436.05 ;
        RECT  66.9 425.4 68.1 426.6 ;
        RECT  51.0 425.4 52.2 426.6 ;
        RECT  70.8 76.8 75.3 78.0 ;
        RECT  74.1 74.1 75.3 75.3 ;
        RECT  72.9 72.6 74.1 75.3 ;
        RECT  69.6 75.0 70.8 78.0 ;
        RECT  60.0 77.1 69.6 78.0 ;
        RECT  65.1 72.6 72.9 73.8 ;
        RECT  61.8 71.7 63.0 74.7 ;
        RECT  58.8 76.8 60.0 78.0 ;
        RECT  59.7 73.5 60.9 74.7 ;
        RECT  58.2 73.5 59.7 74.4 ;
        RECT  57.3 73.5 58.2 75.9 ;
        RECT  51.0 75.0 57.3 75.9 ;
        RECT  56.4 71.7 61.8 72.6 ;
        RECT  55.2 71.7 56.4 73.8 ;
        RECT  52.8 71.7 54.0 73.8 ;
        RECT  49.8 75.0 51.0 76.2 ;
        RECT  45.3 76.8 46.5 78.3 ;
        RECT  33.6 77.4 45.3 78.3 ;
        RECT  43.2 74.1 47.7 75.3 ;
        RECT  42.3 74.1 43.2 76.5 ;
        RECT  35.4 75.6 42.3 76.5 ;
        RECT  40.8 71.7 52.8 72.6 ;
        RECT  39.6 71.7 40.8 73.8 ;
        RECT  36.3 71.7 37.5 74.7 ;
        RECT  34.5 75.0 35.4 76.5 ;
        RECT  32.4 76.8 33.6 78.3 ;
        RECT  33.3 73.5 34.5 75.9 ;
        RECT  24.6 75.0 33.3 75.9 ;
        RECT  30.0 71.7 36.3 72.6 ;
        RECT  28.8 71.7 30.0 73.8 ;
        RECT  26.4 71.7 27.6 73.8 ;
        RECT  23.4 75.0 24.6 76.2 ;
        RECT  17.7 71.7 26.4 72.6 ;
        RECT  16.5 71.7 17.7 75.3 ;
        RECT  15.3 74.1 16.5 75.3 ;
        RECT  15.3 69.0 75.3 70.2 ;
        RECT  70.8 61.2 75.3 62.4 ;
        RECT  74.1 63.9 75.3 65.1 ;
        RECT  72.9 63.9 74.1 66.6 ;
        RECT  69.6 61.2 70.8 64.2 ;
        RECT  60.0 61.2 69.6 62.1 ;
        RECT  65.1 65.4 72.9 66.6 ;
        RECT  61.8 64.5 63.0 67.5 ;
        RECT  58.8 61.2 60.0 62.4 ;
        RECT  59.7 64.5 60.9 65.7 ;
        RECT  58.2 64.8 59.7 65.7 ;
        RECT  57.3 63.3 58.2 65.7 ;
        RECT  51.0 63.3 57.3 64.2 ;
        RECT  56.4 66.6 61.8 67.5 ;
        RECT  55.2 65.4 56.4 67.5 ;
        RECT  52.8 65.4 54.0 67.5 ;
        RECT  49.8 63.0 51.0 64.2 ;
        RECT  45.3 60.9 46.5 62.4 ;
        RECT  33.6 60.9 45.3 61.8 ;
        RECT  43.2 63.9 47.7 65.1 ;
        RECT  42.3 62.7 43.2 65.1 ;
        RECT  35.4 62.7 42.3 63.6 ;
        RECT  40.8 66.6 52.8 67.5 ;
        RECT  39.6 65.4 40.8 67.5 ;
        RECT  36.3 64.5 37.5 67.5 ;
        RECT  34.5 62.7 35.4 64.2 ;
        RECT  32.4 60.9 33.6 62.4 ;
        RECT  33.3 63.3 34.5 65.7 ;
        RECT  24.6 63.3 33.3 64.2 ;
        RECT  30.0 66.6 36.3 67.5 ;
        RECT  28.8 65.4 30.0 67.5 ;
        RECT  26.4 65.4 27.6 67.5 ;
        RECT  23.4 63.0 24.6 64.2 ;
        RECT  17.7 66.6 26.4 67.5 ;
        RECT  16.5 63.9 17.7 67.5 ;
        RECT  15.3 63.9 16.5 65.1 ;
        RECT  15.3 69.0 75.3 70.2 ;
        RECT  70.8 56.4 75.3 57.6 ;
        RECT  74.1 53.7 75.3 54.9 ;
        RECT  72.9 52.2 74.1 54.9 ;
        RECT  69.6 54.6 70.8 57.6 ;
        RECT  60.0 56.7 69.6 57.6 ;
        RECT  65.1 52.2 72.9 53.4 ;
        RECT  61.8 51.3 63.0 54.3 ;
        RECT  58.8 56.4 60.0 57.6 ;
        RECT  59.7 53.1 60.9 54.3 ;
        RECT  58.2 53.1 59.7 54.0 ;
        RECT  57.3 53.1 58.2 55.5 ;
        RECT  51.0 54.6 57.3 55.5 ;
        RECT  56.4 51.3 61.8 52.2 ;
        RECT  55.2 51.3 56.4 53.4 ;
        RECT  52.8 51.3 54.0 53.4 ;
        RECT  49.8 54.6 51.0 55.8 ;
        RECT  45.3 56.4 46.5 57.9 ;
        RECT  33.6 57.0 45.3 57.9 ;
        RECT  43.2 53.7 47.7 54.9 ;
        RECT  42.3 53.7 43.2 56.1 ;
        RECT  35.4 55.2 42.3 56.1 ;
        RECT  40.8 51.3 52.8 52.2 ;
        RECT  39.6 51.3 40.8 53.4 ;
        RECT  36.3 51.3 37.5 54.3 ;
        RECT  34.5 54.6 35.4 56.1 ;
        RECT  32.4 56.4 33.6 57.9 ;
        RECT  33.3 53.1 34.5 55.5 ;
        RECT  24.6 54.6 33.3 55.5 ;
        RECT  30.0 51.3 36.3 52.2 ;
        RECT  28.8 51.3 30.0 53.4 ;
        RECT  26.4 51.3 27.6 53.4 ;
        RECT  23.4 54.6 24.6 55.8 ;
        RECT  17.7 51.3 26.4 52.2 ;
        RECT  16.5 51.3 17.7 54.9 ;
        RECT  15.3 53.7 16.5 54.9 ;
        RECT  15.3 48.6 75.3 49.8 ;
        RECT  70.8 40.8 75.3 42.0 ;
        RECT  74.1 43.5 75.3 44.7 ;
        RECT  72.9 43.5 74.1 46.2 ;
        RECT  69.6 40.8 70.8 43.8 ;
        RECT  60.0 40.8 69.6 41.7 ;
        RECT  65.1 45.0 72.9 46.2 ;
        RECT  61.8 44.1 63.0 47.1 ;
        RECT  58.8 40.8 60.0 42.0 ;
        RECT  59.7 44.1 60.9 45.3 ;
        RECT  58.2 44.4 59.7 45.3 ;
        RECT  57.3 42.9 58.2 45.3 ;
        RECT  51.0 42.9 57.3 43.8 ;
        RECT  56.4 46.2 61.8 47.1 ;
        RECT  55.2 45.0 56.4 47.1 ;
        RECT  52.8 45.0 54.0 47.1 ;
        RECT  49.8 42.6 51.0 43.8 ;
        RECT  45.3 40.5 46.5 42.0 ;
        RECT  33.6 40.5 45.3 41.4 ;
        RECT  43.2 43.5 47.7 44.7 ;
        RECT  42.3 42.3 43.2 44.7 ;
        RECT  35.4 42.3 42.3 43.2 ;
        RECT  40.8 46.2 52.8 47.1 ;
        RECT  39.6 45.0 40.8 47.1 ;
        RECT  36.3 44.1 37.5 47.1 ;
        RECT  34.5 42.3 35.4 43.8 ;
        RECT  32.4 40.5 33.6 42.0 ;
        RECT  33.3 42.9 34.5 45.3 ;
        RECT  24.6 42.9 33.3 43.8 ;
        RECT  30.0 46.2 36.3 47.1 ;
        RECT  28.8 45.0 30.0 47.1 ;
        RECT  26.4 45.0 27.6 47.1 ;
        RECT  23.4 42.6 24.6 43.8 ;
        RECT  17.7 46.2 26.4 47.1 ;
        RECT  16.5 43.5 17.7 47.1 ;
        RECT  15.3 43.5 16.5 44.7 ;
        RECT  15.3 48.6 75.3 49.8 ;
        RECT  128.55 6.0 129.45 6.9 ;
        RECT  124.5 6.0 129.0 6.9 ;
        RECT  128.55 6.45 129.45 12.45 ;
        RECT  124.05 6.0 125.25 7.2 ;
        RECT  138.75 6.0 139.65 6.9 ;
        RECT  134.7 6.0 139.2 6.9 ;
        RECT  138.75 6.45 139.65 12.45 ;
        RECT  134.25 6.0 135.45 7.2 ;
        RECT  148.95 6.0 149.85 6.9 ;
        RECT  144.9 6.0 149.4 6.9 ;
        RECT  148.95 6.45 149.85 12.45 ;
        RECT  144.45 6.0 145.65 7.2 ;
        RECT  128.55 0.3 129.75 1.5 ;
        RECT  138.75 0.3 139.95 1.5 ;
        RECT  148.95 0.3 150.15 1.5 ;
        RECT  90.6 88.8 91.8 90.0 ;
        RECT  90.9 73.5 92.1 74.7 ;
        RECT  72.0 73.5 73.2 74.7 ;
        RECT  87.9 104.7 89.1 105.9 ;
        RECT  88.2 64.8 89.4 66.0 ;
        RECT  72.0 64.8 73.2 66.0 ;
        RECT  85.2 147.6 86.4 148.8 ;
        RECT  85.5 53.1 86.7 54.3 ;
        RECT  72.0 53.1 73.2 54.3 ;
        RECT  82.5 163.5 83.7 164.7 ;
        RECT  82.8 44.4 84.0 45.6 ;
        RECT  72.0 44.4 73.2 45.6 ;
        RECT  114.0 33.3 115.2 34.5 ;
        RECT  108.6 28.65 109.8 29.85 ;
        RECT  111.3 26.25 112.5 27.45 ;
        RECT  114.0 446.4 115.2 447.6 ;
        RECT  116.7 97.95 117.9 99.15 ;
        RECT  119.4 196.05 120.6 197.25 ;
        RECT  16.5 76.5 17.7 77.7 ;
        RECT  16.2 76.8 17.4 78.0 ;
        RECT  106.2 83.1 107.4 84.3 ;
        RECT  105.9 456.6 107.1 457.8 ;
        RECT  95.1 437.1 97.5 438.3 ;
        RECT  133.8 437.1 135.0 438.3 ;
        RECT  144.0 437.1 145.2 438.3 ;
        RECT  154.2 437.1 155.4 438.3 ;
        RECT  122.7 437.1 123.9 438.3 ;
        RECT  101.7 8.1 104.1 9.3 ;
        RECT  133.5 8.1 134.7 9.3 ;
        RECT  133.5 8.1 134.7 9.3 ;
        RECT  153.9 8.1 155.1 9.3 ;
        RECT  87.75 229.05 88.95 230.25 ;
        RECT  87.75 258.45 88.95 259.65 ;
        RECT  87.75 287.85 88.95 289.05 ;
        RECT  87.75 317.25 88.95 318.45 ;
        RECT  87.75 346.65 88.95 347.85 ;
        RECT  87.75 376.05 88.95 377.25 ;
        RECT  87.75 405.45 88.95 406.65 ;
        RECT  87.75 434.85 88.95 436.05 ;
        RECT  95.1 140.55 97.5 141.75 ;
        RECT  95.1 199.35 97.5 200.55 ;
        RECT  75.0 69.15 76.2 70.35 ;
        RECT  95.1 69.15 97.5 70.35 ;
        RECT  75.0 69.15 76.2 70.35 ;
        RECT  95.1 69.15 97.5 70.35 ;
        RECT  75.0 48.75 76.2 49.95 ;
        RECT  95.1 48.75 97.5 49.95 ;
        RECT  75.0 48.75 76.2 49.95 ;
        RECT  95.1 48.75 97.5 49.95 ;
        RECT  -66.3 148.2 -7.5 149.1 ;
        RECT  -66.3 150.9 -7.5 151.8 ;
        RECT  -66.3 153.6 -7.5 154.5 ;
        RECT  -66.3 156.3 -7.5 157.2 ;
        RECT  -66.3 159.0 -7.5 159.9 ;
        RECT  -66.3 161.7 -7.5 162.6 ;
        RECT  -66.3 211.5 -7.5 212.4 ;
        RECT  -66.3 214.2 -7.5 215.1 ;
        RECT  -66.3 216.9 -7.5 217.8 ;
        RECT  -66.3 219.6 -7.5 220.5 ;
        RECT  -56.55 145.5 -55.65 149.1 ;
        RECT  -56.55 145.5 -55.65 149.1 ;
        RECT  -36.15 145.5 -35.25 149.1 ;
        RECT  -7.5 161.7 -3.0 162.6 ;
        RECT  -14.1 88.5 -3.0 89.4 ;
        RECT  -14.7 175.5 -3.0 176.4 ;
        RECT  -7.5 211.5 -3.0 212.4 ;
        RECT  -14.7 180.0 -3.0 180.9 ;
        RECT  -64.5 141.0 -63.3 145.5 ;
        RECT  -61.8 144.3 -60.6 145.5 ;
        RECT  -61.8 143.1 -59.1 144.3 ;
        RECT  -64.5 139.8 -61.5 141.0 ;
        RECT  -64.5 130.2 -63.6 139.8 ;
        RECT  -60.3 135.3 -59.1 143.1 ;
        RECT  -61.2 132.0 -58.2 133.2 ;
        RECT  -64.5 129.0 -63.3 130.2 ;
        RECT  -61.2 129.9 -60.0 131.1 ;
        RECT  -60.9 128.4 -60.0 129.9 ;
        RECT  -62.4 127.5 -60.0 128.4 ;
        RECT  -62.4 121.2 -61.5 127.5 ;
        RECT  -59.1 126.6 -58.2 132.0 ;
        RECT  -60.3 125.4 -58.2 126.6 ;
        RECT  -60.3 123.0 -58.2 124.2 ;
        RECT  -62.7 120.0 -61.5 121.2 ;
        RECT  -64.8 115.5 -63.3 116.7 ;
        RECT  -64.8 103.8 -63.9 115.5 ;
        RECT  -61.8 113.4 -60.6 117.9 ;
        RECT  -63.0 112.5 -60.6 113.4 ;
        RECT  -63.0 105.6 -62.1 112.5 ;
        RECT  -59.1 111.0 -58.2 123.0 ;
        RECT  -60.3 109.8 -58.2 111.0 ;
        RECT  -61.2 106.5 -58.2 107.7 ;
        RECT  -63.0 104.7 -61.5 105.6 ;
        RECT  -64.8 102.6 -63.3 103.8 ;
        RECT  -62.4 103.5 -60.0 104.7 ;
        RECT  -62.4 94.8 -61.5 103.5 ;
        RECT  -59.1 100.2 -58.2 106.5 ;
        RECT  -60.3 99.0 -58.2 100.2 ;
        RECT  -60.3 96.6 -58.2 97.8 ;
        RECT  -62.7 93.6 -61.5 94.8 ;
        RECT  -59.1 87.9 -58.2 96.6 ;
        RECT  -61.8 86.7 -58.2 87.9 ;
        RECT  -61.8 85.5 -60.6 86.7 ;
        RECT  -56.7 85.5 -55.5 145.5 ;
        RECT  -48.9 141.0 -47.7 145.5 ;
        RECT  -51.6 144.3 -50.4 145.5 ;
        RECT  -53.1 143.1 -50.4 144.3 ;
        RECT  -50.7 139.8 -47.7 141.0 ;
        RECT  -48.6 130.2 -47.7 139.8 ;
        RECT  -53.1 135.3 -51.9 143.1 ;
        RECT  -54.0 132.0 -51.0 133.2 ;
        RECT  -48.9 129.0 -47.7 130.2 ;
        RECT  -52.2 129.9 -51.0 131.1 ;
        RECT  -52.2 128.4 -51.3 129.9 ;
        RECT  -52.2 127.5 -49.8 128.4 ;
        RECT  -50.7 121.2 -49.8 127.5 ;
        RECT  -54.0 126.6 -53.1 132.0 ;
        RECT  -54.0 125.4 -51.9 126.6 ;
        RECT  -54.0 123.0 -51.9 124.2 ;
        RECT  -50.7 120.0 -49.5 121.2 ;
        RECT  -48.9 115.5 -47.4 116.7 ;
        RECT  -48.3 103.8 -47.4 115.5 ;
        RECT  -51.6 113.4 -50.4 117.9 ;
        RECT  -51.6 112.5 -49.2 113.4 ;
        RECT  -50.1 105.6 -49.2 112.5 ;
        RECT  -54.0 111.0 -53.1 123.0 ;
        RECT  -54.0 109.8 -51.9 111.0 ;
        RECT  -54.0 106.5 -51.0 107.7 ;
        RECT  -50.7 104.7 -49.2 105.6 ;
        RECT  -48.9 102.6 -47.4 103.8 ;
        RECT  -52.2 103.5 -49.8 104.7 ;
        RECT  -50.7 94.8 -49.8 103.5 ;
        RECT  -54.0 100.2 -53.1 106.5 ;
        RECT  -54.0 99.0 -51.9 100.2 ;
        RECT  -54.0 96.6 -51.9 97.8 ;
        RECT  -50.7 93.6 -49.5 94.8 ;
        RECT  -54.0 87.9 -53.1 96.6 ;
        RECT  -54.0 86.7 -50.4 87.9 ;
        RECT  -51.6 85.5 -50.4 86.7 ;
        RECT  -56.7 85.5 -55.5 145.5 ;
        RECT  -44.1 141.0 -42.9 145.5 ;
        RECT  -41.4 144.3 -40.2 145.5 ;
        RECT  -41.4 143.1 -38.7 144.3 ;
        RECT  -44.1 139.8 -41.1 141.0 ;
        RECT  -44.1 130.2 -43.2 139.8 ;
        RECT  -39.9 135.3 -38.7 143.1 ;
        RECT  -40.8 132.0 -37.8 133.2 ;
        RECT  -44.1 129.0 -42.9 130.2 ;
        RECT  -40.8 129.9 -39.6 131.1 ;
        RECT  -40.5 128.4 -39.6 129.9 ;
        RECT  -42.0 127.5 -39.6 128.4 ;
        RECT  -42.0 121.2 -41.1 127.5 ;
        RECT  -38.7 126.6 -37.8 132.0 ;
        RECT  -39.9 125.4 -37.8 126.6 ;
        RECT  -39.9 123.0 -37.8 124.2 ;
        RECT  -42.3 120.0 -41.1 121.2 ;
        RECT  -44.4 115.5 -42.9 116.7 ;
        RECT  -44.4 103.8 -43.5 115.5 ;
        RECT  -41.4 113.4 -40.2 117.9 ;
        RECT  -42.6 112.5 -40.2 113.4 ;
        RECT  -42.6 105.6 -41.7 112.5 ;
        RECT  -38.7 111.0 -37.8 123.0 ;
        RECT  -39.9 109.8 -37.8 111.0 ;
        RECT  -40.8 106.5 -37.8 107.7 ;
        RECT  -42.6 104.7 -41.1 105.6 ;
        RECT  -44.4 102.6 -42.9 103.8 ;
        RECT  -42.0 103.5 -39.6 104.7 ;
        RECT  -42.0 94.8 -41.1 103.5 ;
        RECT  -38.7 100.2 -37.8 106.5 ;
        RECT  -39.9 99.0 -37.8 100.2 ;
        RECT  -39.9 96.6 -37.8 97.8 ;
        RECT  -42.3 93.6 -41.1 94.8 ;
        RECT  -38.7 87.9 -37.8 96.6 ;
        RECT  -41.4 86.7 -37.8 87.9 ;
        RECT  -41.4 85.5 -40.2 86.7 ;
        RECT  -36.3 85.5 -35.1 145.5 ;
        RECT  -19.65 99.9 -18.45 101.1 ;
        RECT  -14.1 100.05 -13.2 100.95 ;
        RECT  -13.65 100.05 -7.65 100.95 ;
        RECT  -14.25 99.9 -13.05 101.1 ;
        RECT  -19.65 95.1 -18.45 96.3 ;
        RECT  -14.1 95.25 -13.2 96.15 ;
        RECT  -13.65 95.25 -7.65 96.15 ;
        RECT  -14.25 95.1 -13.05 96.3 ;
        RECT  -43.65 236.1 -41.85 237.9 ;
        RECT  -14.85 265.8 -13.65 267.0 ;
        RECT  -14.85 256.2 -13.65 257.4 ;
        RECT  -31.65 247.8 -30.45 249.0 ;
        RECT  -31.65 257.4 -30.45 258.6 ;
        RECT  -14.85 260.4 -13.65 261.6 ;
        RECT  -14.55 257.4 -13.65 261.6 ;
        RECT  -14.85 250.8 -13.65 252.0 ;
        RECT  -14.55 247.5 -13.65 249.0 ;
        RECT  -31.2 247.5 -30.3 249.0 ;
        RECT  -14.55 248.25 -13.65 252.0 ;
        RECT  -31.65 247.8 -30.75 248.25 ;
        RECT  -14.7 247.65 -13.5 248.85 ;
        RECT  -31.35 247.65 -30.15 248.85 ;
        RECT  -31.65 253.2 -30.45 254.4 ;
        RECT  -31.65 253.2 -30.75 257.4 ;
        RECT  -53.55 258.3 -51.75 268.8 ;
        RECT  -55.95 255.3 -54.75 268.8 ;
        RECT  -58.95 255.3 -57.75 268.8 ;
        RECT  -55.95 254.1 -53.25 255.3 ;
        RECT  -58.95 254.1 -57.45 255.3 ;
        RECT  -62.55 254.1 -61.35 268.8 ;
        RECT  -53.55 239.4 -51.15 249.9 ;
        RECT  -55.95 239.4 -54.75 252.9 ;
        RECT  -58.95 239.4 -57.75 252.9 ;
        RECT  -55.95 252.9 -53.25 254.1 ;
        RECT  -58.95 252.9 -57.45 254.1 ;
        RECT  -62.55 239.4 -61.35 254.1 ;
        RECT  -53.55 228.9 -51.15 239.4 ;
        RECT  -55.95 225.9 -54.75 239.4 ;
        RECT  -58.95 225.9 -57.75 239.4 ;
        RECT  -55.95 224.7 -53.25 225.9 ;
        RECT  -58.95 224.7 -57.45 225.9 ;
        RECT  -62.55 224.7 -61.35 239.4 ;
        RECT  -43.05 235.35 -41.85 236.55 ;
        RECT  -32.7 238.05 -31.8 238.95 ;
        RECT  -45.0 238.2 -44.1 239.1 ;
        RECT  -44.55 238.2 -32.25 239.1 ;
        RECT  -32.85 237.9 -31.65 239.1 ;
        RECT  -45.15 238.05 -43.95 239.25 ;
        RECT  -55.8 271.05 -54.9 271.95 ;
        RECT  -55.8 254.1 -54.9 271.65 ;
        RECT  -55.95 270.9 -54.75 272.1 ;
        RECT  -13.65 220.5 -12.75 221.4 ;
        RECT  -32.1 220.65 -31.2 221.55 ;
        RECT  -13.65 221.1 -12.75 241.35 ;
        RECT  -32.1 211.5 -31.2 221.1 ;
        RECT  -13.8 220.35 -12.6 221.55 ;
        RECT  -32.25 220.5 -31.05 221.7 ;
        RECT  -32.85 271.2 -31.65 272.4 ;
        RECT  -13.8 239.55 -12.6 240.75 ;
        RECT  -13.65 251.85 -12.75 252.75 ;
        RECT  -50.1 251.85 -49.2 252.75 ;
        RECT  -13.65 241.35 -12.75 252.3 ;
        RECT  -44.55 251.85 -13.2 252.75 ;
        RECT  -49.65 251.85 -44.55 252.75 ;
        RECT  -50.1 231.3 -49.2 252.3 ;
        RECT  -50.25 249.6 -49.05 250.8 ;
        RECT  -45.9 244.65 -45.0 245.55 ;
        RECT  -45.9 197.55 -45.0 245.1 ;
        RECT  -46.05 244.5 -44.85 245.7 ;
        RECT  -45.9 264.75 -45.0 265.65 ;
        RECT  -45.9 237.75 -45.0 265.2 ;
        RECT  -46.05 264.6 -44.85 265.8 ;
        RECT  -8.4 229.95 -7.5 230.85 ;
        RECT  -8.4 172.2 -7.5 173.1 ;
        RECT  -37.8 172.35 -36.9 173.25 ;
        RECT  -8.4 172.8 -7.5 230.4 ;
        RECT  -37.8 172.8 -36.9 193.8 ;
        RECT  -8.55 229.8 -7.35 231.0 ;
        RECT  -8.55 172.05 -7.35 173.25 ;
        RECT  -37.95 172.2 -36.75 173.4 ;
        RECT  -46.65 292.65 -45.45 293.85 ;
        RECT  -43.2 267.0 -42.3 267.9 ;
        RECT  -43.2 277.5 -42.3 278.4 ;
        RECT  -43.2 267.45 -42.3 278.1 ;
        RECT  -43.35 266.85 -42.15 268.05 ;
        RECT  -43.35 277.35 -42.15 278.55 ;
        RECT  -45.9 316.5 -45.0 317.4 ;
        RECT  -45.9 292.65 -45.0 317.1 ;
        RECT  -46.05 316.35 -44.85 317.55 ;
        RECT  -43.2 267.0 -42.3 267.9 ;
        RECT  -43.2 253.5 -42.3 254.4 ;
        RECT  -43.2 254.1 -42.3 267.45 ;
        RECT  -43.35 266.85 -42.15 268.05 ;
        RECT  -43.35 253.35 -42.15 254.55 ;
        RECT  -45.9 344.7 -45.0 345.6 ;
        RECT  -45.9 292.65 -45.0 345.3 ;
        RECT  -46.05 344.55 -44.85 345.75 ;
        RECT  -62.4 229.95 -61.5 230.85 ;
        RECT  -62.4 177.3 -61.5 230.4 ;
        RECT  -62.55 229.8 -61.35 231.0 ;
        RECT  -52.2 229.95 -51.3 230.85 ;
        RECT  -52.2 177.3 -51.3 230.4 ;
        RECT  -52.35 229.8 -51.15 231.0 ;
        RECT  -25.05 169.8 -23.85 175.8 ;
        RECT  -32.7 165.6 -31.8 171.9 ;
        RECT  -34.5 165.6 -33.6 174.3 ;
        RECT  -33.6 173.1 -31.8 174.3 ;
        RECT  -26.25 169.8 -25.05 171.0 ;
        RECT  -26.25 174.6 -25.05 175.8 ;
        RECT  -33.0 170.7 -31.8 171.9 ;
        RECT  -33.9 165.3 -32.7 166.5 ;
        RECT  -33.0 173.1 -31.8 174.3 ;
        RECT  -36.0 165.3 -34.8 166.5 ;
        RECT  -49.95 169.8 -48.75 175.8 ;
        RECT  -42.0 165.6 -41.1 171.9 ;
        RECT  -40.2 165.6 -39.3 174.3 ;
        RECT  -42.0 173.1 -40.2 174.3 ;
        RECT  -49.95 169.8 -48.75 171.0 ;
        RECT  -49.95 174.6 -48.75 175.8 ;
        RECT  -43.2 170.7 -42.0 171.9 ;
        RECT  -42.3 165.3 -41.1 166.5 ;
        RECT  -43.2 173.1 -42.0 174.3 ;
        RECT  -40.2 165.3 -39.0 166.5 ;
        RECT  -40.8 144.3 -39.6 145.5 ;
        RECT  -40.8 150.9 -39.6 152.1 ;
        RECT  -44.25 144.3 -43.05 145.5 ;
        RECT  -44.25 153.6 -43.05 154.8 ;
        RECT  -64.65 144.3 -63.45 145.5 ;
        RECT  -64.65 156.3 -63.45 157.5 ;
        RECT  -49.05 144.3 -47.85 145.5 ;
        RECT  -49.05 159.0 -47.85 160.2 ;
        RECT  -17.4 153.6 -16.2 154.8 ;
        RECT  -14.1 161.7 -12.9 162.9 ;
        RECT  -27.45 161.7 -26.25 162.9 ;
        RECT  -33.0 153.6 -31.8 154.8 ;
        RECT  -34.8 156.3 -33.6 157.5 ;
        RECT  -47.85 161.7 -46.65 162.9 ;
        RECT  -42.3 159.0 -41.1 160.2 ;
        RECT  -40.5 156.3 -39.3 157.5 ;
        RECT  -16.05 121.05 -15.15 121.95 ;
        RECT  -5.85 121.05 -4.95 121.95 ;
        RECT  -5.7 150.9 -4.8 151.8 ;
        RECT  -15.6 121.05 -5.25 121.95 ;
        RECT  -7.5 150.9 -5.25 151.8 ;
        RECT  -16.2 120.9 -15.0 122.1 ;
        RECT  -6.0 120.9 -4.8 122.1 ;
        RECT  -5.85 150.75 -4.65 151.95 ;
        RECT  -30.9 214.2 -29.7 215.4 ;
        RECT  -44.4 211.5 -43.2 212.7 ;
        RECT  -15.0 216.9 -13.8 218.1 ;
        RECT  -4.05 214.2 -3.15 215.1 ;
        RECT  -7.5 214.2 -3.45 215.1 ;
        RECT  -4.2 214.05 -3.0 215.25 ;
        RECT  -43.35 217.2 -42.15 218.4 ;
        RECT  -43.35 236.4 -42.15 237.6 ;
        RECT  -22.95 219.6 -21.75 220.8 ;
        RECT  -52.35 219.6 -51.15 220.8 ;
        RECT  -8.25 148.2 -7.05 149.4 ;
        RECT  -14.7 126.45 -13.8 127.35 ;
        RECT  -27.75 126.45 -26.85 127.35 ;
        RECT  -27.15 126.45 -14.25 127.35 ;
        RECT  -14.85 126.3 -13.65 127.5 ;
        RECT  -27.9 126.3 -26.7 127.5 ;
        RECT  -27.6 85.5 -26.4 86.7 ;
        RECT  -27.3 85.8 -26.1 87.0 ;
        RECT  -4.5 162.0 -3.3 163.2 ;
        RECT  -14.1 88.5 -12.9 89.7 ;
        RECT  -4.5 88.8 -3.3 90.0 ;
        RECT  -15.0 175.5 -13.8 176.7 ;
        RECT  -4.5 175.8 -3.3 177.0 ;
        RECT  -4.5 211.8 -3.3 213.0 ;
        RECT  -15.0 180.0 -13.8 181.2 ;
        RECT  -4.5 180.3 -3.3 181.5 ;
        RECT  105.3 85.8 106.5 87.0 ;
        RECT  113.4 162.0 114.6 163.2 ;
        RECT  110.7 88.8 111.9 90.0 ;
        RECT  108.0 175.8 109.2 177.0 ;
        RECT  116.1 211.8 117.3 213.0 ;
        RECT  118.8 180.3 120.0 181.5 ;
        RECT  0.0 219.6 2.4 220.8 ;
        RECT  95.4 230.7 98.1 231.9 ;
        RECT  -8.1 230.7 -6.9 231.9 ;
        Layer  via2 ; 
        RECT  125.1 152.7 125.7 153.3 ;
        RECT  135.3 152.7 135.9 153.3 ;
        RECT  145.5 152.7 146.1 153.3 ;
        RECT  128.7 32.4 129.3 33.0 ;
        RECT  138.9 32.4 139.5 33.0 ;
        RECT  149.1 32.4 149.7 33.0 ;
        RECT  128.7 32.7 129.3 33.3 ;
        RECT  138.9 32.7 139.5 33.3 ;
        RECT  149.1 32.7 149.7 33.3 ;
        RECT  16.8 74.4 17.4 75.0 ;
        RECT  16.8 64.2 17.4 64.8 ;
        RECT  16.8 54.0 17.4 54.6 ;
        RECT  16.8 43.8 17.4 44.4 ;
        RECT  124.35 6.3 124.95 6.9 ;
        RECT  134.55 6.3 135.15 6.9 ;
        RECT  144.75 6.3 145.35 6.9 ;
        RECT  128.85 0.6 129.45 1.2 ;
        RECT  139.05 0.6 139.65 1.2 ;
        RECT  149.25 0.6 149.85 1.2 ;
        RECT  91.2 73.8 91.8 74.4 ;
        RECT  72.3 73.8 72.9 74.4 ;
        RECT  88.5 65.1 89.1 65.7 ;
        RECT  72.3 65.1 72.9 65.7 ;
        RECT  85.8 53.4 86.4 54.0 ;
        RECT  72.3 53.4 72.9 54.0 ;
        RECT  83.1 44.7 83.7 45.3 ;
        RECT  72.3 44.7 72.9 45.3 ;
        RECT  16.5 77.1 17.1 77.7 ;
        RECT  106.5 83.4 107.1 84.0 ;
        RECT  -61.5 87.0 -60.9 87.6 ;
        RECT  -51.3 87.0 -50.7 87.6 ;
        RECT  -41.1 87.0 -40.5 87.6 ;
        RECT  -14.4 247.95 -13.8 248.55 ;
        RECT  -31.05 247.95 -30.45 248.55 ;
        RECT  -43.05 217.5 -42.45 218.1 ;
        RECT  -43.05 236.7 -42.45 237.3 ;
        RECT  -27.0 86.1 -26.4 86.7 ;
        RECT  -4.2 162.3 -3.6 162.9 ;
        RECT  -4.2 89.1 -3.6 89.7 ;
        RECT  -4.2 176.1 -3.6 176.7 ;
        RECT  -4.2 212.1 -3.6 212.7 ;
        RECT  -4.2 180.6 -3.6 181.2 ;
        RECT  105.6 86.1 106.2 86.7 ;
        RECT  113.7 162.3 114.3 162.9 ;
        RECT  111.0 89.1 111.6 89.7 ;
        RECT  108.3 176.1 108.9 176.7 ;
        RECT  116.4 212.1 117.0 212.7 ;
        RECT  119.1 180.6 119.7 181.2 ;
        RECT  95.7 231.0 96.3 231.6 ;
        RECT  97.2 231.0 97.8 231.6 ;
        RECT  -7.8 231.0 -7.2 231.6 ;
        Layer  metal3 ; 
        RECT  -27.15 85.5 105.9 87.0 ;
        RECT  -3.0 161.7 114.0 163.2 ;
        RECT  -3.0 88.5 111.3 90.0 ;
        RECT  -3.0 175.5 108.6 177.0 ;
        RECT  -3.0 211.5 116.7 213.0 ;
        RECT  -3.0 180.0 119.4 181.5 ;
        RECT  -6.6 230.4 95.1 231.9 ;
        RECT  128.25 0.0 129.75 30.15 ;
        RECT  138.45 0.0 139.95 30.15 ;
        RECT  148.65 0.0 150.15 30.15 ;
        RECT  73.5 73.2 91.5 74.7 ;
        RECT  73.5 64.5 88.8 66.0 ;
        RECT  73.5 52.8 86.1 54.3 ;
        RECT  73.5 44.1 83.4 45.6 ;
        RECT  0.0 73.95 17.1 75.45 ;
        RECT  0.0 63.75 17.1 65.25 ;
        RECT  0.0 53.55 17.1 55.05 ;
        RECT  0.0 43.35 17.1 44.85 ;
        RECT  124.5 152.1 126.3 153.9 ;
        RECT  134.7 152.1 136.5 153.9 ;
        RECT  144.9 152.1 146.7 153.9 ;
        RECT  128.1 31.8 129.9 33.6 ;
        RECT  138.3 31.8 140.1 33.6 ;
        RECT  148.5 31.8 150.3 33.6 ;
        RECT  128.1 32.1 129.9 33.9 ;
        RECT  138.3 32.1 140.1 33.9 ;
        RECT  148.5 32.1 150.3 33.9 ;
        RECT  16.2 73.8 18.0 75.6 ;
        RECT  16.2 63.6 18.0 65.4 ;
        RECT  16.2 53.4 18.0 55.2 ;
        RECT  16.2 43.2 18.0 45.0 ;
        RECT  123.75 153.75 125.25 155.25 ;
        RECT  123.75 6.45 125.25 154.5 ;
        RECT  124.5 153.75 126.15 155.25 ;
        RECT  123.75 5.7 125.55 7.5 ;
        RECT  133.95 153.75 135.45 155.25 ;
        RECT  133.95 6.45 135.45 154.5 ;
        RECT  134.7 153.75 136.35 155.25 ;
        RECT  133.95 5.7 135.75 7.5 ;
        RECT  144.15 153.75 145.65 155.25 ;
        RECT  144.15 6.45 145.65 154.5 ;
        RECT  144.9 153.75 146.55 155.25 ;
        RECT  144.15 5.7 145.95 7.5 ;
        RECT  128.25 0.0 130.05 1.8 ;
        RECT  138.45 0.0 140.25 1.8 ;
        RECT  148.65 0.0 150.45 1.8 ;
        RECT  90.6 73.2 92.4 75.0 ;
        RECT  71.7 73.2 73.5 75.0 ;
        RECT  87.9 64.5 89.7 66.3 ;
        RECT  71.7 64.5 73.5 66.3 ;
        RECT  85.2 52.8 87.0 54.6 ;
        RECT  71.7 52.8 73.5 54.6 ;
        RECT  82.5 44.1 84.3 45.9 ;
        RECT  71.7 44.1 73.5 45.9 ;
        RECT  15.9 76.5 17.7 78.3 ;
        RECT  16.95 82.8 18.45 84.3 ;
        RECT  16.95 76.5 18.45 83.55 ;
        RECT  17.7 82.8 106.2 84.3 ;
        RECT  105.9 82.8 107.7 84.6 ;
        RECT  -43.35 216.9 -41.85 236.55 ;
        RECT  -62.1 86.4 -60.3 88.2 ;
        RECT  -51.9 86.4 -50.1 88.2 ;
        RECT  -41.7 86.4 -39.9 88.2 ;
        RECT  -14.55 247.5 -13.65 249.0 ;
        RECT  -31.2 247.5 -30.3 249.0 ;
        RECT  -31.2 247.5 -14.1 249.0 ;
        RECT  -15.0 247.35 -13.2 249.15 ;
        RECT  -31.65 247.35 -29.85 249.15 ;
        RECT  -43.65 216.9 -41.85 218.7 ;
        RECT  -43.65 236.1 -41.85 237.9 ;
        RECT  -27.6 85.5 -25.8 87.3 ;
        RECT  -4.8 161.7 -3.0 163.5 ;
        RECT  -4.8 88.5 -3.0 90.3 ;
        RECT  -4.8 175.5 -3.0 177.3 ;
        RECT  -4.8 211.5 -3.0 213.3 ;
        RECT  -4.8 180.0 -3.0 181.8 ;
        RECT  105.0 85.5 106.8 87.3 ;
        RECT  113.1 161.7 114.9 163.5 ;
        RECT  110.4 88.5 112.2 90.3 ;
        RECT  107.7 175.5 109.5 177.3 ;
        RECT  115.8 211.5 117.6 213.3 ;
        RECT  118.5 180.0 120.3 181.8 ;
        RECT  95.1 230.4 98.4 232.2 ;
        RECT  -8.4 230.4 -6.6 232.2 ;
    END 
END    ecc 
END    LIBRARY 
